magic
tech sky130A
timestamp 1717366634
<< pwell >>
rect -760 -150 760 150
<< nnmos >>
rect -646 -21 -596 21
rect -508 -21 -458 21
rect -370 -21 -320 21
rect -232 -21 -182 21
rect -94 -21 -44 21
rect 44 -21 94 21
rect 182 -21 232 21
rect 320 -21 370 21
rect 458 -21 508 21
rect 596 -21 646 21
<< mvndiff >>
rect -675 15 -646 21
rect -675 -15 -669 15
rect -652 -15 -646 15
rect -675 -21 -646 -15
rect -596 15 -567 21
rect -596 -15 -590 15
rect -573 -15 -567 15
rect -596 -21 -567 -15
rect -537 15 -508 21
rect -537 -15 -531 15
rect -514 -15 -508 15
rect -537 -21 -508 -15
rect -458 15 -429 21
rect -458 -15 -452 15
rect -435 -15 -429 15
rect -458 -21 -429 -15
rect -399 15 -370 21
rect -399 -15 -393 15
rect -376 -15 -370 15
rect -399 -21 -370 -15
rect -320 15 -291 21
rect -320 -15 -314 15
rect -297 -15 -291 15
rect -320 -21 -291 -15
rect -261 15 -232 21
rect -261 -15 -255 15
rect -238 -15 -232 15
rect -261 -21 -232 -15
rect -182 15 -153 21
rect -182 -15 -176 15
rect -159 -15 -153 15
rect -182 -21 -153 -15
rect -123 15 -94 21
rect -123 -15 -117 15
rect -100 -15 -94 15
rect -123 -21 -94 -15
rect -44 15 -15 21
rect -44 -15 -38 15
rect -21 -15 -15 15
rect -44 -21 -15 -15
rect 15 15 44 21
rect 15 -15 21 15
rect 38 -15 44 15
rect 15 -21 44 -15
rect 94 15 123 21
rect 94 -15 100 15
rect 117 -15 123 15
rect 94 -21 123 -15
rect 153 15 182 21
rect 153 -15 159 15
rect 176 -15 182 15
rect 153 -21 182 -15
rect 232 15 261 21
rect 232 -15 238 15
rect 255 -15 261 15
rect 232 -21 261 -15
rect 291 15 320 21
rect 291 -15 297 15
rect 314 -15 320 15
rect 291 -21 320 -15
rect 370 15 399 21
rect 370 -15 376 15
rect 393 -15 399 15
rect 370 -21 399 -15
rect 429 15 458 21
rect 429 -15 435 15
rect 452 -15 458 15
rect 429 -21 458 -15
rect 508 15 537 21
rect 508 -15 514 15
rect 531 -15 537 15
rect 508 -21 537 -15
rect 567 15 596 21
rect 567 -15 573 15
rect 590 -15 596 15
rect 567 -21 596 -15
rect 646 15 675 21
rect 646 -15 652 15
rect 669 -15 675 15
rect 646 -21 675 -15
<< mvndiffc >>
rect -669 -15 -652 15
rect -590 -15 -573 15
rect -531 -15 -514 15
rect -452 -15 -435 15
rect -393 -15 -376 15
rect -314 -15 -297 15
rect -255 -15 -238 15
rect -176 -15 -159 15
rect -117 -15 -100 15
rect -38 -15 -21 15
rect 21 -15 38 15
rect 100 -15 117 15
rect 159 -15 176 15
rect 238 -15 255 15
rect 297 -15 314 15
rect 376 -15 393 15
rect 435 -15 452 15
rect 514 -15 531 15
rect 573 -15 590 15
rect 652 -15 669 15
<< mvpsubdiff >>
rect -742 103 742 132
rect -742 -103 -713 103
rect 713 78 742 103
rect 713 -78 719 78
rect 736 -78 742 78
rect 713 -103 742 -78
rect -742 -132 742 -103
<< mvpsubdiffcont >>
rect 719 -78 736 78
<< poly >>
rect -646 57 -596 65
rect -646 40 -638 57
rect -604 40 -596 57
rect -646 21 -596 40
rect -508 57 -458 65
rect -508 40 -500 57
rect -466 40 -458 57
rect -508 21 -458 40
rect -370 57 -320 65
rect -370 40 -362 57
rect -328 40 -320 57
rect -370 21 -320 40
rect -232 57 -182 65
rect -232 40 -224 57
rect -190 40 -182 57
rect -232 21 -182 40
rect -94 57 -44 65
rect -94 40 -86 57
rect -52 40 -44 57
rect -94 21 -44 40
rect 44 57 94 65
rect 44 40 52 57
rect 86 40 94 57
rect 44 21 94 40
rect 182 57 232 65
rect 182 40 190 57
rect 224 40 232 57
rect 182 21 232 40
rect 320 57 370 65
rect 320 40 328 57
rect 362 40 370 57
rect 320 21 370 40
rect 458 57 508 65
rect 458 40 466 57
rect 500 40 508 57
rect 458 21 508 40
rect 596 57 646 65
rect 596 40 604 57
rect 638 40 646 57
rect 596 21 646 40
rect -646 -40 -596 -21
rect -646 -57 -638 -40
rect -604 -57 -596 -40
rect -646 -65 -596 -57
rect -508 -40 -458 -21
rect -508 -57 -500 -40
rect -466 -57 -458 -40
rect -508 -65 -458 -57
rect -370 -40 -320 -21
rect -370 -57 -362 -40
rect -328 -57 -320 -40
rect -370 -65 -320 -57
rect -232 -40 -182 -21
rect -232 -57 -224 -40
rect -190 -57 -182 -40
rect -232 -65 -182 -57
rect -94 -40 -44 -21
rect -94 -57 -86 -40
rect -52 -57 -44 -40
rect -94 -65 -44 -57
rect 44 -40 94 -21
rect 44 -57 52 -40
rect 86 -57 94 -40
rect 44 -65 94 -57
rect 182 -40 232 -21
rect 182 -57 190 -40
rect 224 -57 232 -40
rect 182 -65 232 -57
rect 320 -40 370 -21
rect 320 -57 328 -40
rect 362 -57 370 -40
rect 320 -65 370 -57
rect 458 -40 508 -21
rect 458 -57 466 -40
rect 500 -57 508 -40
rect 458 -65 508 -57
rect 596 -40 646 -21
rect 596 -57 604 -40
rect 638 -57 646 -40
rect 596 -65 646 -57
<< polycont >>
rect -638 40 -604 57
rect -500 40 -466 57
rect -362 40 -328 57
rect -224 40 -190 57
rect -86 40 -52 57
rect 52 40 86 57
rect 190 40 224 57
rect 328 40 362 57
rect 466 40 500 57
rect 604 40 638 57
rect -638 -57 -604 -40
rect -500 -57 -466 -40
rect -362 -57 -328 -40
rect -224 -57 -190 -40
rect -86 -57 -52 -40
rect 52 -57 86 -40
rect 190 -57 224 -40
rect 328 -57 362 -40
rect 466 -57 500 -40
rect 604 -57 638 -40
<< locali >>
rect 719 78 736 86
rect -646 40 -638 57
rect -604 40 -596 57
rect -508 40 -500 57
rect -466 40 -458 57
rect -370 40 -362 57
rect -328 40 -320 57
rect -232 40 -224 57
rect -190 40 -182 57
rect -94 40 -86 57
rect -52 40 -44 57
rect 44 40 52 57
rect 86 40 94 57
rect 182 40 190 57
rect 224 40 232 57
rect 320 40 328 57
rect 362 40 370 57
rect 458 40 466 57
rect 500 40 508 57
rect 596 40 604 57
rect 638 40 646 57
rect -669 15 -652 23
rect -669 -23 -652 -15
rect -590 15 -573 23
rect -590 -23 -573 -15
rect -531 15 -514 23
rect -531 -23 -514 -15
rect -452 15 -435 23
rect -452 -23 -435 -15
rect -393 15 -376 23
rect -393 -23 -376 -15
rect -314 15 -297 23
rect -314 -23 -297 -15
rect -255 15 -238 23
rect -255 -23 -238 -15
rect -176 15 -159 23
rect -176 -23 -159 -15
rect -117 15 -100 23
rect -117 -23 -100 -15
rect -38 15 -21 23
rect -38 -23 -21 -15
rect 21 15 38 23
rect 21 -23 38 -15
rect 100 15 117 23
rect 100 -23 117 -15
rect 159 15 176 23
rect 159 -23 176 -15
rect 238 15 255 23
rect 238 -23 255 -15
rect 297 15 314 23
rect 297 -23 314 -15
rect 376 15 393 23
rect 376 -23 393 -15
rect 435 15 452 23
rect 435 -23 452 -15
rect 514 15 531 23
rect 514 -23 531 -15
rect 573 15 590 23
rect 573 -23 590 -15
rect 652 15 669 23
rect 652 -23 669 -15
rect -646 -57 -638 -40
rect -604 -57 -596 -40
rect -508 -57 -500 -40
rect -466 -57 -458 -40
rect -370 -57 -362 -40
rect -328 -57 -320 -40
rect -232 -57 -224 -40
rect -190 -57 -182 -40
rect -94 -57 -86 -40
rect -52 -57 -44 -40
rect 44 -57 52 -40
rect 86 -57 94 -40
rect 182 -57 190 -40
rect 224 -57 232 -40
rect 320 -57 328 -40
rect 362 -57 370 -40
rect 458 -57 466 -40
rect 500 -57 508 -40
rect 596 -57 604 -40
rect 638 -57 646 -40
rect 719 -86 736 -78
<< viali >>
rect -638 40 -604 57
rect -500 40 -466 57
rect -362 40 -328 57
rect -224 40 -190 57
rect -86 40 -52 57
rect 52 40 86 57
rect 190 40 224 57
rect 328 40 362 57
rect 466 40 500 57
rect 604 40 638 57
rect -669 -15 -652 15
rect -590 -15 -573 15
rect -531 -15 -514 15
rect -452 -15 -435 15
rect -393 -15 -376 15
rect -314 -15 -297 15
rect -255 -15 -238 15
rect -176 -15 -159 15
rect -117 -15 -100 15
rect -38 -15 -21 15
rect 21 -15 38 15
rect 100 -15 117 15
rect 159 -15 176 15
rect 238 -15 255 15
rect 297 -15 314 15
rect 376 -15 393 15
rect 435 -15 452 15
rect 514 -15 531 15
rect 573 -15 590 15
rect 652 -15 669 15
rect -638 -57 -604 -40
rect -500 -57 -466 -40
rect -362 -57 -328 -40
rect -224 -57 -190 -40
rect -86 -57 -52 -40
rect 52 -57 86 -40
rect 190 -57 224 -40
rect 328 -57 362 -40
rect 466 -57 500 -40
rect 604 -57 638 -40
<< metal1 >>
rect -644 57 -598 60
rect -644 40 -638 57
rect -604 40 -598 57
rect -644 37 -598 40
rect -506 57 -460 60
rect -506 40 -500 57
rect -466 40 -460 57
rect -506 37 -460 40
rect -368 57 -322 60
rect -368 40 -362 57
rect -328 40 -322 57
rect -368 37 -322 40
rect -230 57 -184 60
rect -230 40 -224 57
rect -190 40 -184 57
rect -230 37 -184 40
rect -92 57 -46 60
rect -92 40 -86 57
rect -52 40 -46 57
rect -92 37 -46 40
rect 46 57 92 60
rect 46 40 52 57
rect 86 40 92 57
rect 46 37 92 40
rect 184 57 230 60
rect 184 40 190 57
rect 224 40 230 57
rect 184 37 230 40
rect 322 57 368 60
rect 322 40 328 57
rect 362 40 368 57
rect 322 37 368 40
rect 460 57 506 60
rect 460 40 466 57
rect 500 40 506 57
rect 460 37 506 40
rect 598 57 644 60
rect 598 40 604 57
rect 638 40 644 57
rect 598 37 644 40
rect -672 15 -649 21
rect -672 -15 -669 15
rect -652 -15 -649 15
rect -672 -21 -649 -15
rect -593 15 -570 21
rect -593 -15 -590 15
rect -573 -15 -570 15
rect -593 -21 -570 -15
rect -534 15 -511 21
rect -534 -15 -531 15
rect -514 -15 -511 15
rect -534 -21 -511 -15
rect -455 15 -432 21
rect -455 -15 -452 15
rect -435 -15 -432 15
rect -455 -21 -432 -15
rect -396 15 -373 21
rect -396 -15 -393 15
rect -376 -15 -373 15
rect -396 -21 -373 -15
rect -317 15 -294 21
rect -317 -15 -314 15
rect -297 -15 -294 15
rect -317 -21 -294 -15
rect -258 15 -235 21
rect -258 -15 -255 15
rect -238 -15 -235 15
rect -258 -21 -235 -15
rect -179 15 -156 21
rect -179 -15 -176 15
rect -159 -15 -156 15
rect -179 -21 -156 -15
rect -120 15 -97 21
rect -120 -15 -117 15
rect -100 -15 -97 15
rect -120 -21 -97 -15
rect -41 15 -18 21
rect -41 -15 -38 15
rect -21 -15 -18 15
rect -41 -21 -18 -15
rect 18 15 41 21
rect 18 -15 21 15
rect 38 -15 41 15
rect 18 -21 41 -15
rect 97 15 120 21
rect 97 -15 100 15
rect 117 -15 120 15
rect 97 -21 120 -15
rect 156 15 179 21
rect 156 -15 159 15
rect 176 -15 179 15
rect 156 -21 179 -15
rect 235 15 258 21
rect 235 -15 238 15
rect 255 -15 258 15
rect 235 -21 258 -15
rect 294 15 317 21
rect 294 -15 297 15
rect 314 -15 317 15
rect 294 -21 317 -15
rect 373 15 396 21
rect 373 -15 376 15
rect 393 -15 396 15
rect 373 -21 396 -15
rect 432 15 455 21
rect 432 -15 435 15
rect 452 -15 455 15
rect 432 -21 455 -15
rect 511 15 534 21
rect 511 -15 514 15
rect 531 -15 534 15
rect 511 -21 534 -15
rect 570 15 593 21
rect 570 -15 573 15
rect 590 -15 593 15
rect 570 -21 593 -15
rect 649 15 672 21
rect 649 -15 652 15
rect 669 -15 672 15
rect 649 -21 672 -15
rect -644 -40 -598 -37
rect -644 -57 -638 -40
rect -604 -57 -598 -40
rect -644 -60 -598 -57
rect -506 -40 -460 -37
rect -506 -57 -500 -40
rect -466 -57 -460 -40
rect -506 -60 -460 -57
rect -368 -40 -322 -37
rect -368 -57 -362 -40
rect -328 -57 -322 -40
rect -368 -60 -322 -57
rect -230 -40 -184 -37
rect -230 -57 -224 -40
rect -190 -57 -184 -40
rect -230 -60 -184 -57
rect -92 -40 -46 -37
rect -92 -57 -86 -40
rect -52 -57 -46 -40
rect -92 -60 -46 -57
rect 46 -40 92 -37
rect 46 -57 52 -40
rect 86 -57 92 -40
rect 46 -60 92 -57
rect 184 -40 230 -37
rect 184 -57 190 -40
rect 224 -57 230 -40
rect 184 -60 230 -57
rect 322 -40 368 -37
rect 322 -57 328 -40
rect 362 -57 368 -40
rect 322 -60 368 -57
rect 460 -40 506 -37
rect 460 -57 466 -40
rect 500 -57 506 -40
rect 460 -60 506 -57
rect 598 -40 644 -37
rect 598 -57 604 -40
rect 638 -57 644 -40
rect 598 -60 644 -57
<< properties >>
string FIXED_BBOX -727 -117 727 117
string gencell sky130_fd_pr__nfet_03v3_nvt
string library sky130
string parameters w 0.42 l 0.5 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 0 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
