* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_R72FWE a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt GSense_nFET_10VD_5Vg_1nf VD_H VG_H VLow_Src VSUBS
XXM1 VLow_Src VSUBS VD_H VG_H sky130_fd_pr__nfet_g5v0d10v5_R72FWE
.ends

.subckt GSense_Contacts_nFT_g5_10Vd_1nf VSUBS
XGSense_nFET_10VD_5Vg_1nf_0 GSense_nFET_10VD_5Vg_1nf_0/VD_H GSense_nFET_10VD_5Vg_1nf_0/VG_H
+ GSense_nFET_10VD_5Vg_1nf_0/VLow_Src VSUBS GSense_nFET_10VD_5Vg_1nf
.ends

.subckt sky130_fd_pr__nfet_01v8_J36GRF a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt GSense_nFET_1f1WL150n_V1 VD_H VG_H VLow_Src VSUBS
XXM3 VD_H VG_H VLow_Src VSUBS sky130_fd_pr__nfet_01v8_J36GRF
.ends

.subckt GSense_nFET_1W015L_1F_Contacts GSense_nFET_1f1WL150n_V1_0/VG_H VSUBS
XGSense_nFET_1f1WL150n_V1_0 GSense_nFET_1f1WL150n_V1_0/VD_H GSense_nFET_1f1WL150n_V1_0/VG_H
+ GSense_nFET_1f1WL150n_V1_0/VLow_Src VSUBS GSense_nFET_1f1WL150n_V1
.ends

.subckt sky130_fd_pr__nfet_03v3_nvt_XW2EXC a_n4524_n42# a_3638_n42# a_n3538_n42# a_n1764_n42#
+ a_5746_n130# a_n3914_n130# a_n3638_n130# a_6240_n42# a_n778_n42# a_2100_n42# a_50_n42#
+ a_3480_n42# a_n6950_n130# a_878_n42# a_n6674_n130# a_n5352_n42# a_n6398_n130# a_n4366_n42#
+ a_n1212_n42# a_4466_n42# a_n1982_n130# a_n2592_n42# a_3814_n130# a_3538_n130# a_n4800_n42#
+ a_n226_n42# a_n3814_n42# a_3914_n42# a_n1706_n130# a_326_n42# a_6850_n130# a_2928_n42#
+ a_n6180_n42# a_6574_n130# a_n4742_n130# a_n5194_n42# a_n2040_n42# a_5294_n42# a_6298_n130#
+ a_1882_n130# a_1154_n42# a_n1054_n42# a_n4466_n130# a_6516_n42# a_n4642_n42# a_4742_n42#
+ a_1606_n130# a_1982_n42# a_3756_n42# a_n1882_n42# a_168_n42# a_502_n130# a_n5628_n42#
+ a_4642_n130# a_n2868_n42# a_n502_n42# a_226_n130# a_602_n42# a_4366_n130# a_n2810_n130#
+ a_n2534_n130# a_996_n42# a_5570_n42# a_n2258_n130# a_n5470_n42# a_3204_n42# a_n1330_n42#
+ a_1430_n42# a_4584_n42# a_n602_n130# a_n5570_n130# a_n326_n130# a_n6456_n42# a_n5294_n130#
+ a_n3696_n42# a_n2316_n42# a_2710_n130# a_444_n42# a_2434_n130# a_n5904_n42# a_n5018_n130#
+ a_2158_n130# a_n4918_n42# a_4032_n42# a_5470_n130# a_1272_n42# a_5018_n42# a_5194_n130#
+ a_n3144_n42# a_6398_n42# a_n6298_n42# a_2258_n42# a_n3362_n130# a_n2158_n42# a_4860_n42#
+ a_n3086_n130# a_n6732_n42# a_n5746_n42# a_n384_n42# a_5846_n42# a_n3972_n42# a_n1606_n42#
+ a_1706_n42# a_n2986_n42# a_720_n42# a_n6122_n130# a_3086_n42# a_3262_n130# a_n1430_n130#
+ a_n1154_n130# a_n3420_n42# a_6674_n42# a_n6574_n42# a_4308_n42# a_n2434_n42# a_2534_n42#
+ a_5688_n42# a_1548_n42# a_n4190_n130# a_n660_n42# a_6022_n130# a_1330_n130# a_6122_n42#
+ a_1054_n130# a_778_n130# a_n6022_n42# a_5136_n42# a_n3262_n42# a_3362_n42# a_2376_n42#
+ a_n7008_n42# a_4090_n130# a_4918_n130# a_n4248_n42# a_6950_n42# a_n6850_n42# a_n2710_n42#
+ a_n1488_n42# a_2810_n42# a_5964_n42# a_n878_n130# a_1824_n42# a_n108_n42# a_n4090_n42#
+ a_4190_n42# a_n5846_n130# a_2986_n130# a_n50_n130# a_n5076_n42# a_n936_n42# a_5412_n42#
+ a_6792_n42# a_2652_n42# a_n7142_n264# m1_n6988_n248#
X0 a_n6022_n42# a_n6122_n130# a_n6180_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1 a_n3538_n42# a_n3638_n130# a_n3696_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X2 a_3086_n42# a_2986_n130# a_2928_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X3 a_6950_n42# a_6850_n130# a_6792_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X4 a_n3262_n42# a_n3362_n130# a_n3420_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X5 a_5294_n42# a_5194_n130# a_5136_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X6 a_6674_n42# a_6574_n130# a_6516_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X7 a_n4642_n42# a_n4742_n130# a_n4800_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X8 a_n2986_n42# a_n3086_n130# a_n3144_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X9 a_1706_n42# a_1606_n130# a_1548_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X10 a_6398_n42# a_6298_n130# a_6240_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X11 a_n4366_n42# a_n4466_n130# a_n4524_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X12 a_n1882_n42# a_n1982_n130# a_n2040_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X13 a_n502_n42# a_n602_n130# a_n660_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X14 a_1430_n42# a_1330_n130# a_1272_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X15 a_50_n42# a_n50_n130# a_n108_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X16 a_n5746_n42# a_n5846_n130# a_n5904_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X17 a_2810_n42# a_2710_n130# a_2652_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X18 a_n4090_n42# a_n4190_n130# a_n4248_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X19 a_878_n42# a_778_n130# a_720_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X20 a_1154_n42# a_1054_n130# a_996_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X21 a_n226_n42# a_n326_n130# a_n384_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X22 a_n5470_n42# a_n5570_n130# a_n5628_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X23 a_2534_n42# a_2434_n130# a_2376_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X24 a_n5194_n42# a_n5294_n130# a_n5352_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X25 a_n6850_n42# a_n6950_n130# a_n7008_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X26 a_2258_n42# a_2158_n130# a_2100_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X27 a_3914_n42# a_3814_n130# a_3756_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X28 a_6122_n42# a_6022_n130# a_5964_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X29 a_n6574_n42# a_n6674_n130# a_n6732_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X30 a_3638_n42# a_3538_n130# a_3480_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X31 a_n1606_n42# a_n1706_n130# a_n1764_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X32 a_n6298_n42# a_n6398_n130# a_n6456_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X33 a_3362_n42# a_3262_n130# a_3204_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X34 a_5018_n42# a_4918_n130# a_4860_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X35 a_602_n42# a_502_n130# a_444_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X36 a_n1330_n42# a_n1430_n130# a_n1488_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X37 a_4742_n42# a_4642_n130# a_4584_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X38 a_n2710_n42# a_n2810_n130# a_n2868_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X39 a_n1054_n42# a_n1154_n130# a_n1212_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X40 a_326_n42# a_226_n130# a_168_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X41 a_1982_n42# a_1882_n130# a_1824_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X42 a_4466_n42# a_4366_n130# a_4308_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X43 a_n4918_n42# a_n5018_n130# a_n5076_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X44 a_n2434_n42# a_n2534_n130# a_n2592_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X45 a_4190_n42# a_4090_n130# a_4032_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X46 a_5846_n42# a_5746_n130# a_5688_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X47 a_n3814_n42# a_n3914_n130# a_n3972_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X48 a_n2158_n42# a_n2258_n130# a_n2316_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X49 a_n778_n42# a_n878_n130# a_n936_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X50 a_5570_n42# a_5470_n130# a_5412_n42# a_n7142_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
.ends

.subckt GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH VG_H VD_H VLow_Src li_174_n490# VSUBS
XXM1 VLow_Src VD_H VLow_Src VLow_Src VG_H VG_H VG_H VLow_Src VD_H VD_H VLow_Src VLow_Src
+ li_174_n490# VD_H VG_H VD_H VG_H VD_H VLow_Src VLow_Src VG_H VD_H VG_H VG_H VD_H
+ VD_H VD_H VLow_Src VG_H VD_H VG_H VLow_Src VLow_Src VG_H VG_H VLow_Src VD_H VD_H
+ VG_H VG_H VLow_Src VD_H VG_H VD_H VLow_Src VD_H VG_H VD_H VD_H VLow_Src VLow_Src
+ VG_H VLow_Src VG_H VLow_Src VLow_Src VG_H VLow_Src VG_H VG_H VG_H VD_H VLow_Src
+ VG_H VD_H VD_H VLow_Src VD_H VLow_Src VG_H VG_H VG_H VD_H VG_H VD_H VLow_Src VG_H
+ VD_H VG_H VD_H VG_H VG_H VD_H VLow_Src VG_H VLow_Src VLow_Src VG_H VD_H VD_H VLow_Src
+ VLow_Src VG_H VD_H VD_H VG_H VLow_Src VLow_Src VLow_Src VD_H VLow_Src VD_H VLow_Src
+ VLow_Src VLow_Src VG_H VD_H VG_H VG_H VG_H VLow_Src VLow_Src VD_H VD_H VLow_Src
+ VD_H VLow_Src VD_H VG_H VD_H VG_H VG_H VLow_Src VG_H VG_H VD_H VLow_Src VD_H VLow_Src
+ VLow_Src VD_H VG_H VG_H VD_H VD_H VLow_Src VD_H VD_H VLow_Src VD_H VG_H VLow_Src
+ VD_H VLow_Src VD_H VG_H VG_H VG_H VLow_Src VLow_Src VD_H VLow_Src VD_H VSUBS VD_H
+ sky130_fd_pr__nfet_03v3_nvt_XW2EXC
.ends

.subckt nFET_3p3Vd_3VG_51NF_LTherm_Contacts m1_5996_2684# VSUBS
XGSense_nFET_3VD_3Vg_51nf_V2AllGates_VH_0 GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH_0/VG_H
+ GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH_0/VD_H GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH_0/VLow_Src
+ m1_n4654_560# VSUBS GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH
.ends

.subckt GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline VG_H VD_H VLow_Src m1_6800_n480#
+ VSUBS
XXM1 VLow_Src VD_H VLow_Src VLow_Src VG_H VG_H VG_H VLow_Src VD_H VD_H VLow_Src VLow_Src
+ VG_H VD_H VG_H VD_H VG_H VD_H VLow_Src VLow_Src VG_H VD_H VG_H VG_H VD_H VD_H VD_H
+ VLow_Src VG_H VD_H VG_H VLow_Src VLow_Src VG_H VG_H VLow_Src VD_H VD_H VG_H VG_H
+ VLow_Src VD_H VG_H VD_H VLow_Src VD_H VG_H VD_H VD_H VLow_Src VLow_Src VG_H VLow_Src
+ VG_H VLow_Src VLow_Src VG_H VLow_Src VG_H VG_H VG_H VD_H VLow_Src VG_H VD_H VD_H
+ VLow_Src VD_H VLow_Src VG_H VG_H m1_6800_n480# VD_H VG_H VD_H VLow_Src VG_H VD_H
+ VG_H VD_H VG_H VG_H VD_H VLow_Src VG_H VLow_Src VLow_Src VG_H VD_H VD_H VLow_Src
+ VLow_Src VG_H VD_H VD_H VG_H VLow_Src VLow_Src VLow_Src VD_H VLow_Src VD_H VLow_Src
+ VLow_Src VLow_Src VG_H VD_H VG_H VG_H VG_H VLow_Src VLow_Src VD_H VD_H VLow_Src
+ VD_H VLow_Src VD_H VG_H VD_H VG_H VG_H VLow_Src VG_H VG_H VD_H VLow_Src VD_H VLow_Src
+ VLow_Src VD_H VG_H VG_H VD_H VD_H VLow_Src VD_H VD_H VLow_Src VD_H VG_H VLow_Src
+ VD_H VLow_Src VD_H VG_H VG_H VG_H VLow_Src VLow_Src VD_H VLow_Src VD_H VSUBS VD_H
+ sky130_fd_pr__nfet_03v3_nvt_XW2EXC
.ends

.subckt nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts m1_5996_6595# VSUBS
XGSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0 GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0/VG_H
+ GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0/VD_H GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0/VLow_Src
+ m2_n1290_6370# VSUBS GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_W5U4AW c2_n3079_n3000# m4_n3179_n3100#
X0 c2_n3079_n3000# m4_n3179_n3100# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
.ends

.subckt sky130_fd_sc_hvl__buf_8 VPWR VPB VNB VGND X A
X0 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5 M=8
X1 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5 M=8
X2 a_45_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.2025 ps=1.29 w=0.75 l=0.5 M=3
X3 VPWR A a_45_443# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5 M=3
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ a_n683_n200# a_n189_n297# a_29_n297# a_189_n200#
+ a_n901_n200# a_247_n297# a_n407_n297# a_465_n297# a_407_n200# a_n625_n297# a_683_n297#
+ a_625_n200# a_n843_n297# w_n1101_n497# a_843_n200# a_n29_n200# a_n247_n200# a_n465_n200#
X0 a_n247_n200# a_n407_n297# a_n465_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X1 a_843_n200# a_683_n297# a_625_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X2 a_407_n200# a_247_n297# a_189_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X3 a_189_n200# a_29_n297# a_n29_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X4 a_n465_n200# a_n625_n297# a_n683_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X5 a_625_n200# a_465_n297# a_407_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X6 a_n29_n200# a_n189_n297# a_n247_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X7 a_n683_n200# a_n843_n297# a_n901_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_TGFUGS a_n792_n200# a_298_n200# a_516_n200# a_734_n200#
+ a_n926_n422# a_138_n288# a_n298_n288# a_80_n200# a_356_n288# a_n516_n288# a_574_n288#
+ a_n734_n288# a_n138_n200# a_n356_n200# a_n574_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X1 a_n574_n200# a_n734_n288# a_n792_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
X2 a_734_n200# a_574_n288# a_516_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X3 a_298_n200# a_138_n288# a_80_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X4 a_n138_n200# a_n298_n288# a_n356_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X5 a_n356_n200# a_n516_n288# a_n574_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X6 a_516_n200# a_356_n288# a_298_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_S5N9F3 a_124_2496# a_n4122_n2932# a_n4122_2496#
+ a_2054_n2932# a_2054_2496# a_896_n2932# a_510_2496# a_3598_2496# a_3984_2496# a_3598_n2932#
+ a_2440_2496# a_n3736_n2932# a_1668_n2932# a_n1806_n2932# a_5142_n2932# a_510_n2932#
+ a_n2192_2496# a_n3736_2496# a_3212_n2932# a_n5410_n3062# a_1668_2496# a_n262_2496#
+ a_4756_n2932# a_5142_2496# a_2826_n2932# a_n2192_n2932# a_n1806_2496# a_n5280_2496#
+ a_n648_n2932# a_n5280_n2932# a_n3350_n2932# a_4756_2496# a_3212_2496# a_1282_n2932#
+ a_124_n2932# a_n1420_n2932# a_n4894_n2932# a_896_2496# a_n2964_n2932# a_n3350_2496#
+ a_n4508_2496# a_n4894_2496# a_n4508_n2932# a_4370_n2932# a_1282_2496# a_2826_2496#
+ a_2440_n2932# a_3984_n2932# a_n1034_2496# a_n2578_2496# a_n1420_2496# a_n2964_2496#
+ a_n262_n2932# a_n648_2496# a_n1034_n2932# a_4370_2496# a_n2578_n2932#
X0 a_n262_2496# a_n262_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X1 a_n3350_2496# a_n3350_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X2 a_n4122_2496# a_n4122_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X3 a_n4894_2496# a_n4894_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X4 a_n3736_2496# a_n3736_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X5 a_1282_2496# a_1282_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X6 a_5142_2496# a_5142_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X7 a_4756_2496# a_4756_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X8 a_124_2496# a_124_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X9 a_510_2496# a_510_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X10 a_896_2496# a_896_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X11 a_n5280_2496# a_n5280_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X12 a_n648_2496# a_n648_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X13 a_n4508_2496# a_n4508_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X14 a_n2192_2496# a_n2192_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X15 a_n1034_2496# a_n1034_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X16 a_2054_2496# a_2054_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X17 a_1668_2496# a_1668_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X18 a_2440_2496# a_2440_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X19 a_n1420_2496# a_n1420_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X20 a_n2578_2496# a_n2578_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X21 a_n1806_2496# a_n1806_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X22 a_3212_2496# a_3212_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X23 a_3598_2496# a_3598_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X24 a_n2964_2496# a_n2964_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X25 a_4370_2496# a_4370_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X26 a_2826_2496# a_2826_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X27 a_3984_2496# a_3984_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_3YBPVB a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_sc_hvl__schmittbuf_1 X A VPB VNB VPWR VGND
X0 X a_117_181# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.315925 ps=1.45 w=0.75 l=0.5
X1 a_217_207# a_117_181# a_64_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.5
X2 VPWR A a_231_463# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.34075 pd=1.73 as=0.105 ps=1.03 w=0.75 l=0.5
X3 VGND A a_217_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.315925 pd=1.45 as=0.0588 ps=0.7 w=0.42 l=0.5
X4 a_78_463# VGND VNB sky130_fd_pr__res_generic_nd__hv w=0.29 l=1.355
X5 a_64_207# VPWR VPB sky130_fd_pr__res_generic_pd__hv w=0.29 l=3.11
X6 X a_117_181# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.34075 ps=1.73 w=1.5 l=0.5
X7 a_231_463# A a_117_181# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X8 a_231_463# a_117_181# a_78_463# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X9 a_217_207# A a_117_181# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YUHPXE a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PKVMTM a_80_n200# a_n272_n422# a_n138_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n272_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC a_80_n200# a_n272_n422# a_n138_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n272_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_WRT4AW c1_n3036_n3000# m3_n3136_n3100#
X0 c1_n3036_n3000# m3_n3136_n3100# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YEUEBV a_n792_n200# a_138_n297# a_n298_n297#
+ a_298_n200# a_356_n297# a_n516_n297# a_574_n297# a_516_n200# a_n734_n297# a_734_n200#
+ a_n80_n297# a_80_n200# a_n138_n200# a_n356_n200# a_n574_n200# w_n992_n497#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X1 a_n574_n200# a_n734_n297# a_n792_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
X2 a_734_n200# a_574_n297# a_516_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X3 a_298_n200# a_138_n297# a_80_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X4 a_n138_n200# a_n298_n297# a_n356_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X5 a_n356_n200# a_n516_n297# a_n574_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X6 a_516_n200# a_356_n297# a_298_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YUHPBG a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_sc_hvl__inv_8 VNB VGND VPWR VPB Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5 M=8
X1 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.1575 pd=1.17 as=0.105 ps=1.03 w=0.75 l=0.5 M=8
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__fill_4 abstract view
.subckt sky130_fd_sc_hvl__fill_4 VNB VGND VPWR VPB
.ends

.subckt example_por vdd3v3 vdd1v8 vss porb_h por_l porb_l
Xsky130_fd_pr__cap_mim_m3_2_W5U4AW_0 vss sky130_fd_sc_hvl__schmittbuf_1_0/A sky130_fd_pr__cap_mim_m3_2_W5U4AW
Xsky130_fd_sc_hvl__buf_8_1 vdd1v8 vdd1v8 vss vss porb_l sky130_fd_sc_hvl__inv_8_0/A
+ sky130_fd_sc_hvl__buf_8
Xsky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ_0 m1_502_7653# m1_502_7653# m1_502_7653# m1_502_7653#
+ vdd3v3 m1_502_7653# m1_502_7653# m1_502_7653# vdd3v3 m1_502_7653# m1_502_7653# m1_502_7653#
+ m1_502_7653# vdd3v3 vdd3v3 vdd3v3 m1_502_7653# vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ
Xsky130_fd_pr__nfet_g5v0d10v5_TGFUGS_0 m1_721_6815# vss m1_721_6815# vss vss m1_721_6815#
+ m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# vss
+ m1_721_6815# vss m1_721_6815# sky130_fd_pr__nfet_g5v0d10v5_TGFUGS
Xsky130_fd_pr__res_xhigh_po_0p69_S5N9F3_0 li_5638_5813# li_1391_165# li_1006_5813#
+ li_7567_165# li_7182_5813# li_6023_165# li_5638_5813# li_8726_5813# li_9498_5813#
+ li_9111_165# li_7954_5813# li_1391_165# li_6795_165# li_3707_165# vss li_6023_165#
+ li_3322_5813# li_1778_5813# li_8339_165# vss li_7182_5813# li_4866_5813# li_9883_165#
+ vss li_8339_165# li_2935_165# li_3322_5813# vss li_4479_165# vss li_2163_165# vdd3v3
+ li_8726_5813# li_6795_165# li_5251_165# li_3707_165# li_619_165# li_6410_5813# li_2163_165#
+ li_1778_5813# li_1006_5813# vss li_619_165# li_9883_165# li_6410_5813# li_7954_5813#
+ li_7567_165# li_9111_165# li_4094_5813# li_2550_5813# li_4094_5813# li_2550_5813#
+ li_5251_165# li_4866_5813# li_4479_165# li_9498_5813# li_2935_165# sky130_fd_pr__res_xhigh_po_0p69_S5N9F3
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_0 m1_2756_6573# sky130_fd_sc_hvl__schmittbuf_1_0/A
+ vdd3v3 m1_6249_7690# sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_sc_hvl__schmittbuf_1_0 sky130_fd_sc_hvl__inv_8_0/A sky130_fd_sc_hvl__schmittbuf_1_0/A
+ vdd3v3 vss vdd3v3 vss sky130_fd_sc_hvl__schmittbuf_1
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_1 m1_185_6573# m1_721_6815# vdd3v3 m1_2993_7658#
+ sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_2 m1_2756_6573# m1_4283_8081# vdd3v3 m1_2756_6573#
+ sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_3 m1_185_6573# m1_502_7653# vdd3v3 m1_185_6573#
+ sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_pr__pfet_g5v0d10v5_YUHPXE_0 m1_4283_8081# m1_6249_7690# vdd3v3 vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_YUHPXE
Xsky130_fd_pr__nfet_g5v0d10v5_PKVMTM_0 m1_2756_6573# vss vss m1_721_6815# sky130_fd_pr__nfet_g5v0d10v5_PKVMTM
Xsky130_fd_pr__nfet_g5v0d10v5_ZK8HQC_0 m1_185_6573# vss vss li_2550_5813# sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC
Xsky130_fd_pr__cap_mim_m3_1_WRT4AW_0 sky130_fd_sc_hvl__schmittbuf_1_0/A vss sky130_fd_pr__cap_mim_m3_1_WRT4AW
Xsky130_fd_pr__pfet_g5v0d10v5_YEUEBV_0 vdd3v3 m1_4283_8081# m1_4283_8081# m1_4283_8081#
+ m1_4283_8081# m1_4283_8081# m1_4283_8081# vdd3v3 m1_4283_8081# m1_4283_8081# m1_4283_8081#
+ vdd3v3 m1_4283_8081# vdd3v3 m1_4283_8081# vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_YEUEBV
Xsky130_fd_pr__pfet_g5v0d10v5_YUHPBG_0 m1_502_7653# m1_2993_7658# vdd3v3 vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_YUHPBG
Xsky130_fd_sc_hvl__inv_8_0 vss vss vdd1v8 vdd1v8 por_l sky130_fd_sc_hvl__inv_8_0/A
+ sky130_fd_sc_hvl__inv_8
Xsky130_fd_sc_hvl__fill_4_0 vss vss vdd3v3 vdd3v3 sky130_fd_sc_hvl__fill_4
Xsky130_fd_sc_hvl__buf_8_0 vdd3v3 vdd3v3 vss vss porb_h sky130_fd_sc_hvl__inv_8_0/A
+ sky130_fd_sc_hvl__buf_8
.ends

.subckt user_analog_proj_example example_por_0/por_l example_por_1/por_l example_por_0/vdd1v8
+ example_por_1/vdd3v3 example_por_1/porb_l example_por_0/vdd3v3 example_por_1/porb_h
+ example_por_0/porb_l example_por_0/porb_h VSUBS example_por_1/vdd1v8
Xexample_por_0 example_por_0/vdd3v3 example_por_0/vdd1v8 VSUBS example_por_0/porb_h
+ example_por_0/por_l example_por_0/porb_l example_por
Xexample_por_1 example_por_1/vdd3v3 example_por_1/vdd1v8 VSUBS example_por_1/porb_h
+ example_por_1/por_l example_por_1/porb_l example_por
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_WLCVX2 a_n50_n197# a_50_n100# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n308_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt GSense_pFET_10VD_5Vg_1nf VD_H VLow_Src VG_H
XXM1 VG_H VLow_Src VD_H sky130_fd_pr__pfet_g5v0d10v5_WLCVX2
.ends

.subckt GSense_pFET_10Vd_5p5Vg_1nf
XGSense_pFET_10VD_5Vg_1nf_0 GSense_pFET_10VD_5Vg_1nf_0/VD_H GSense_pFET_10VD_5Vg_1nf_0/VLow_Src
+ GSense_pFET_10VD_5Vg_1nf_0/VG_H GSense_pFET_10VD_5Vg_1nf
.ends

.subckt sky130_fd_pr__nfet_03v3_nvt_J2JJF2 a_858_n42# a_30_n42# a_306_n42# a_n798_n42#
+ a_n1292_n130# a_1134_n42# a_n1016_n130# a_n246_n42# a_1192_n130# a_n1074_n42# a_916_n130#
+ a_n1484_n264# a_188_n42# a_n522_n42# a_n1350_n42# a_n88_n42# a_464_n42# a_n364_n42#
+ a_1292_n42# a_n1192_n42# a_n640_n42# a_740_n42# a_582_n42# a_640_n130# a_364_n130#
+ a_88_n130# a_n740_n130# a_1016_n42# a_n916_n42# a_n188_n130# a_n464_n130#
X0 a_740_n42# a_640_n130# a_582_n42# a_n1484_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1 a_n1192_n42# a_n1292_n130# a_n1350_n42# a_n1484_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X2 a_464_n42# a_364_n130# a_306_n42# a_n1484_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X3 a_n916_n42# a_n1016_n130# a_n1074_n42# a_n1484_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X4 a_188_n42# a_88_n130# a_30_n42# a_n1484_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X5 a_n640_n42# a_n740_n130# a_n798_n42# a_n1484_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X6 a_1292_n42# a_1192_n130# a_1134_n42# a_n1484_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X7 a_n364_n42# a_n464_n130# a_n522_n42# a_n1484_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X8 a_n88_n42# a_n188_n130# a_n246_n42# a_n1484_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X9 a_1016_n42# a_916_n130# a_858_n42# a_n1484_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
.ends

.subckt GSense_nFET_3VD_3Vg_10nf_V2 VG_H VD_H VLow_Src m1_1152_n620# VSUBS
XXM1 VD_H VLow_Src VD_H VD_H VG_H VLow_Src VG_H VD_H VG_H VLow_Src VG_H VSUBS VD_H
+ VLow_Src VD_H VLow_Src VLow_Src VD_H VD_H VLow_Src VLow_Src VD_H VLow_Src VG_H VG_H
+ VG_H VG_H VLow_Src VD_H m1_1152_n620# VG_H sky130_fd_pr__nfet_03v3_nvt_J2JJF2
.ends

.subckt nFET_3VD_3VG_10nF_Contacts m1_5996_2684# VSUBS
XGSense_nFET_3VD_3Vg_10nf_V2_0 GSense_nFET_3VD_3Vg_10nf_V2_0/VG_H GSense_nFET_3VD_3Vg_10nf_V2_0/VD_H
+ GSense_nFET_3VD_3Vg_10nf_V2_0/VLow_Src m1_n1260_1140# VSUBS GSense_nFET_3VD_3Vg_10nf_V2
.ends

.subckt sky130_fd_pr__nfet_03v3_nvt_EJ4KLV a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_03v3_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt GSense_nFET_3VD_3Vg_1nf VD_H VG_H VLow_Src VSUBS
XXM1 VLow_Src VSUBS VD_H VG_H sky130_fd_pr__nfet_03v3_nvt_EJ4KLV
.ends

.subckt GSense_Contacts_nFET_3V_1nf VSUBS
XGSense_nFET_3VD_3Vg_1nf_0 GSense_nFET_3VD_3Vg_1nf_0/VD_H GSense_nFET_3VD_3Vg_1nf_0/VG_H
+ GSense_nFET_3VD_3Vg_1nf_0/VLow_Src VSUBS GSense_nFET_3VD_3Vg_1nf
.ends

.subckt nFET_3VD_3VG_50nF_Therm_FET12 m1_5996_2973# VSUBS
XGSense_nFET_3VD_3Vg_51nf_V2AllGates_Mid_Therm_0 GSense_nFET_3VD_3Vg_51nf_V2AllGates_Mid_Therm_0/VG_H
+ GSense_nFET_3VD_3Vg_51nf_V2AllGates_Mid_Therm_0/VD_H GSense_nFET_3VD_3Vg_51nf_V2AllGates_Mid_Therm_0/VLow_Src
+ m2_n1312_3142# VSUBS GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline
.ends

.subckt sky130_fd_pr__nfet_03v3_nvt_VB5P9F a_50_n42# a_326_n42# a_n226_n42# a_168_n42#
+ a_502_n130# a_602_n42# a_n502_n42# a_226_n130# a_n602_n130# a_n326_n130# a_444_n42#
+ a_n794_n264# a_n384_n42# a_n660_n42# a_n108_n42# a_n50_n130#
X0 a_n502_n42# a_n602_n130# a_n660_n42# a_n794_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1 a_50_n42# a_n50_n130# a_n108_n42# a_n794_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X2 a_n226_n42# a_n326_n130# a_n384_n42# a_n794_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X3 a_602_n42# a_502_n130# a_444_n42# a_n794_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X4 a_326_n42# a_226_n130# a_168_n42# a_n794_n264# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
.ends

.subckt GSense_nFET_3VD_3Vg_5nf_V2 VD_H VG_H VLow_Src m1_672_n216# VSUBS
Xsky130_fd_pr__nfet_03v3_nvt_VB5P9F_0 VLow_Src VD_H VD_H VLow_Src VG_H VLow_Src VLow_Src
+ VG_H VG_H VG_H VD_H VSUBS VLow_Src VD_H VD_H m1_672_n216# sky130_fd_pr__nfet_03v3_nvt_VB5P9F
.ends

.subckt GSense_nFET_3p3V_5nF_Contacts_V2 VSUBS
XGSense_nFET_3VD_3Vg_5nf_V2_1 GSense_nFET_3VD_3Vg_5nf_V2_1/VD_H GSense_nFET_3VD_3Vg_5nf_V2_1/VG_H
+ GSense_nFET_3VD_3Vg_5nf_V2_1/VLow_Src m1_n1260_1140# VSUBS GSense_nFET_3VD_3Vg_5nf_V2
.ends

.subckt sky130_fd_pr__pfet_01v8_8JS3FC a_n73_n100# a_15_n100# a_n33_n197#
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt GSense_pFET_1p8VD_1p8Vg_1nf VD_H VLow_Src VG_H
XXM1 VD_H VLow_Src VG_H sky130_fd_pr__pfet_01v8_8JS3FC
.ends

.subckt GSense_Contacts_pfet_1p8Vd_1p8Vg
XGSense_pFET_1p8VD_1p8Vg_1nf_0 GSense_pFET_1p8VD_1p8Vg_1nf_0/VD_H GSense_pFET_1p8VD_1p8Vg_1nf_0/VLow_Src
+ GSense_pFET_1p8VD_1p8Vg_1nf_0/VG_H GSense_pFET_1p8VD_1p8Vg_1nf
.ends

.subckt user_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11] gpio_analog[12]
+ gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16] gpio_analog[17]
+ gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5] gpio_analog[6]
+ gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10] gpio_noesd[11]
+ gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16] gpio_noesd[17]
+ gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5] gpio_noesd[6]
+ gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10] io_analog[1]
+ io_analog[2] io_analog[3] io_analog[4] io_analog[5] io_analog[6] io_analog[7] io_analog[8]
+ io_analog[9] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i io_analog[4]_uq0 io_analog[4]_uq1 io_analog[4]_uq2 io_analog[4]_uq3
+ io_analog[5]_uq0 io_analog[5]_uq1 io_analog[5]_uq2 io_analog[5]_uq3 io_analog[5]_uq4
+ io_analog[6]_uq0 io_analog[6]_uq1 io_analog[6]_uq2 io_analog[6]_uq3 io_analog[6]_uq4
+ vssa1_uq0 vssa1_uq1 vssd2_uq0 vdda2_uq0 vdda1_uq0 vssd1_uq0 vssa2_uq0 vccd2_uq0
+ vdda1_uq1 vssd1
XGSense_Contacts_nFT_g5_10Vd_1nf_1 vssa1_uq1 GSense_Contacts_nFT_g5_10Vd_1nf
XGSense_Contacts_nFT_g5_10Vd_1nf_2 vssa1_uq1 GSense_Contacts_nFT_g5_10Vd_1nf
XGSense_nFET_1W015L_1F_Contacts_0 GSense_nFET_1W015L_1F_Contacts_0/GSense_nFET_1f1WL150n_V1_0/VG_H
+ vssa1_uq1 GSense_nFET_1W015L_1F_Contacts
XGSense_nFET_1W015L_1F_Contacts_2 GSense_nFET_1W015L_1F_Contacts_2/GSense_nFET_1f1WL150n_V1_0/VG_H
+ vssa1_uq1 GSense_nFET_1W015L_1F_Contacts
XGSense_nFET_1W015L_1F_Contacts_1 GSense_nFET_1W015L_1F_Contacts_1/GSense_nFET_1f1WL150n_V1_0/VG_H
+ vssa1_uq1 GSense_nFET_1W015L_1F_Contacts
XGSense_nFET_1W015L_1F_Contacts_3 GSense_nFET_1W015L_1F_Contacts_3/GSense_nFET_1f1WL150n_V1_0/VG_H
+ vssa1_uq1 GSense_nFET_1W015L_1F_Contacts
XnFET_3p3Vd_3VG_51NF_LTherm_Contacts_0 nFET_3p3Vd_3VG_51NF_LTherm_Contacts_0/m1_5996_2684#
+ vssa1_uq1 nFET_3p3Vd_3VG_51NF_LTherm_Contacts
XnFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_0 nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_0/m1_5996_6595#
+ vssa1_uq1 nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts
XnFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_1 nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_1/m1_5996_6595#
+ vssa1_uq1 nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts
XnFET_3p3Vd_3VG_51NF_LTherm_Contacts_1 gpio_analog[7] vssa1_uq1 nFET_3p3Vd_3VG_51NF_LTherm_Contacts
XGSense_nFET_1W015L_1F_Contacts_4 GSense_nFET_1W015L_1F_Contacts_4/GSense_nFET_1f1WL150n_V1_0/VG_H
+ vssa1_uq1 GSense_nFET_1W015L_1F_Contacts
Xuser_analog_proj_example_0 io_out[16] io_out[12] vccd1 vdda1_uq1 io_out[11] io_analog[4]_uq3
+ gpio_analog[3] io_out[15] gpio_analog[7] vssa1_uq1 vccd1 user_analog_proj_example
XnFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_2 nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_2/m1_5996_6595#
+ vssa1_uq1 nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts
XnFET_3p3Vd_3VG_51NF_LTherm_Contacts_2 nFET_3p3Vd_3VG_51NF_LTherm_Contacts_2/m1_5996_2684#
+ vssa1_uq1 nFET_3p3Vd_3VG_51NF_LTherm_Contacts
XGSense_nFET_1W015L_1F_Contacts_5 GSense_nFET_1W015L_1F_Contacts_5/GSense_nFET_1f1WL150n_V1_0/VG_H
+ vssa1_uq1 GSense_nFET_1W015L_1F_Contacts
XnFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_3 gpio_analog[7] vssa1_uq1 nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts
XnFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_5 nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_5/m1_5996_6595#
+ vssa1_uq1 nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts
XGSense_pFET_10Vd_5p5Vg_1nf_0 GSense_pFET_10Vd_5p5Vg_1nf
XGSense_pFET_10Vd_5p5Vg_1nf_1 GSense_pFET_10Vd_5p5Vg_1nf
XGSense_pFET_10Vd_5p5Vg_1nf_2 GSense_pFET_10Vd_5p5Vg_1nf
XnFET_3VD_3VG_10nF_Contacts_0 nFET_3VD_3VG_10nF_Contacts_0/m1_5996_2684# vssa1_uq1
+ nFET_3VD_3VG_10nF_Contacts
XGSense_Contacts_nFET_3V_1nf_0 vssa1_uq1 GSense_Contacts_nFET_3V_1nf
XnFET_3VD_3VG_10nF_Contacts_1 nFET_3VD_3VG_10nF_Contacts_1/m1_5996_2684# vssa1_uq1
+ nFET_3VD_3VG_10nF_Contacts
XGSense_Contacts_nFET_3V_1nf_1 vssa1_uq1 GSense_Contacts_nFET_3V_1nf
XnFET_3VD_3VG_10nF_Contacts_2 nFET_3VD_3VG_10nF_Contacts_2/m1_5996_2684# vssa1_uq1
+ nFET_3VD_3VG_10nF_Contacts
XnFET_3VD_3VG_50nF_Therm_FET12_0 nFET_3VD_3VG_50nF_Therm_FET12_0/m1_5996_2973# vssa1_uq1
+ nFET_3VD_3VG_50nF_Therm_FET12
XnFET_3VD_3VG_10nF_Contacts_3 gpio_analog[7] vssa1_uq1 nFET_3VD_3VG_10nF_Contacts
XGSense_Contacts_nFET_3V_1nf_2 vssa1_uq1 GSense_Contacts_nFET_3V_1nf
XnFET_3VD_3VG_50nF_Therm_FET12_1 gpio_analog[7] vssa1_uq1 nFET_3VD_3VG_50nF_Therm_FET12
XGSense_Contacts_nFET_3V_1nf_3 vssa1_uq1 GSense_Contacts_nFET_3V_1nf
XGSense_nFET_3p3V_5nF_Contacts_V2_0 vssa1_uq1 GSense_nFET_3p3V_5nF_Contacts_V2
XGSense_Contacts_pfet_1p8Vd_1p8Vg_0 GSense_Contacts_pfet_1p8Vd_1p8Vg
XnFET_3VD_3VG_50nF_Therm_FET12_3 nFET_3VD_3VG_50nF_Therm_FET12_3/m1_5996_2973# vssa1_uq1
+ nFET_3VD_3VG_50nF_Therm_FET12
XGSense_nFET_3p3V_5nF_Contacts_V2_1 vssa1_uq1 GSense_nFET_3p3V_5nF_Contacts_V2
XGSense_Contacts_pfet_1p8Vd_1p8Vg_1 GSense_Contacts_pfet_1p8Vd_1p8Vg
XGSense_nFET_3p3V_5nF_Contacts_V2_2 vssa1_uq1 GSense_nFET_3p3V_5nF_Contacts_V2
XGSense_Contacts_pfet_1p8Vd_1p8Vg_2 GSense_Contacts_pfet_1p8Vd_1p8Vg
XGSense_Contacts_nFT_g5_10Vd_1nf_0 vssa1_uq1 GSense_Contacts_nFT_g5_10Vd_1nf
R0 io_oeb[15] vssd1 sky130_fd_pr__res_generic_m3 w=0.56 l=0.6
R1 io_clamp_high[0] io_analog[4]_uq3 sky130_fd_pr__res_generic_m3 w=11 l=0.25
R2 vssd1 io_oeb[11] sky130_fd_pr__res_generic_m3 w=0.56 l=0.58
R3 io_clamp_low[1] vssa1_uq1 sky130_fd_pr__res_generic_m3 w=11 l=0.25
R4 io_oeb[16] vssd1 sky130_fd_pr__res_generic_m3 w=0.56 l=0.31
R5 io_clamp_low[0] vssa1_uq1 sky130_fd_pr__res_generic_m3 w=11 l=0.25
R6 vssd1 io_oeb[12] sky130_fd_pr__res_generic_m3 w=0.56 l=0.49
R7 io_clamp_high[2] vssa1_uq1 sky130_fd_pr__res_generic_m3 w=11 l=0.25
R8 io_clamp_high[1] vssa1_uq1 sky130_fd_pr__res_generic_m3 w=11 l=0.25
R9 io_clamp_low[2] vssa1_uq1 sky130_fd_pr__res_generic_m3 w=11 l=0.25
.ends

