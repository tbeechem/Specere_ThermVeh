magic
tech sky130A
magscale 1 2
timestamp 1717279825
<< error_p >>
rect -125 114 -67 120
rect 67 114 125 120
rect -125 80 -113 114
rect 67 80 79 114
rect -125 74 -67 80
rect 67 74 125 80
rect -221 -80 -163 -74
rect -29 -80 29 -74
rect 163 -80 221 -74
rect -221 -114 -209 -80
rect -29 -114 -17 -80
rect 163 -114 175 -80
rect -221 -120 -163 -114
rect -29 -120 29 -114
rect 163 -120 221 -114
<< pwell >>
rect -407 -252 407 252
<< nmos >>
rect -207 -42 -177 42
rect -111 -42 -81 42
rect -15 -42 15 42
rect 81 -42 111 42
rect 177 -42 207 42
<< ndiff >>
rect -269 30 -207 42
rect -269 -30 -257 30
rect -223 -30 -207 30
rect -269 -42 -207 -30
rect -177 30 -111 42
rect -177 -30 -161 30
rect -127 -30 -111 30
rect -177 -42 -111 -30
rect -81 30 -15 42
rect -81 -30 -65 30
rect -31 -30 -15 30
rect -81 -42 -15 -30
rect 15 30 81 42
rect 15 -30 31 30
rect 65 -30 81 30
rect 15 -42 81 -30
rect 111 30 177 42
rect 111 -30 127 30
rect 161 -30 177 30
rect 111 -42 177 -30
rect 207 30 269 42
rect 207 -30 223 30
rect 257 -30 269 30
rect 207 -42 269 -30
<< ndiffc >>
rect -257 -30 -223 30
rect -161 -30 -127 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 127 -30 161 30
rect 223 -30 257 30
<< psubdiff >>
rect -371 182 -275 216
rect 275 182 371 216
rect -371 120 -337 182
rect 337 120 371 182
rect -371 -182 -337 -120
rect 337 -182 371 -120
rect -371 -216 -275 -182
rect 275 -216 371 -182
<< psubdiffcont >>
rect -275 182 275 216
rect -371 -120 -337 120
rect 337 -120 371 120
rect -275 -216 275 -182
<< poly >>
rect -129 114 -63 130
rect -129 80 -113 114
rect -79 80 -63 114
rect -207 42 -177 68
rect -129 64 -63 80
rect 63 114 129 130
rect 63 80 79 114
rect 113 80 129 114
rect -111 42 -81 64
rect -15 42 15 68
rect 63 64 129 80
rect 81 42 111 64
rect 177 42 207 68
rect -207 -64 -177 -42
rect -225 -80 -159 -64
rect -111 -68 -81 -42
rect -15 -64 15 -42
rect -225 -114 -209 -80
rect -175 -114 -159 -80
rect -225 -130 -159 -114
rect -33 -80 33 -64
rect 81 -68 111 -42
rect 177 -64 207 -42
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect -33 -130 33 -114
rect 159 -80 225 -64
rect 159 -114 175 -80
rect 209 -114 225 -80
rect 159 -130 225 -114
<< polycont >>
rect -113 80 -79 114
rect 79 80 113 114
rect -209 -114 -175 -80
rect -17 -114 17 -80
rect 175 -114 209 -80
<< locali >>
rect -371 182 -275 216
rect 275 182 371 216
rect -371 120 -337 182
rect 337 120 371 182
rect -129 80 -113 114
rect -79 80 -63 114
rect 63 80 79 114
rect 113 80 129 114
rect -257 30 -223 46
rect -257 -46 -223 -30
rect -161 30 -127 46
rect -161 -46 -127 -30
rect -65 30 -31 46
rect -65 -46 -31 -30
rect 31 30 65 46
rect 31 -46 65 -30
rect 127 30 161 46
rect 127 -46 161 -30
rect 223 30 257 46
rect 223 -46 257 -30
rect -225 -114 -209 -80
rect -175 -114 -159 -80
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect 159 -114 175 -80
rect 209 -114 225 -80
rect -371 -182 -337 -120
rect 337 -182 371 -120
rect -371 -216 -275 -182
rect 275 -216 371 -182
<< viali >>
rect -113 80 -79 114
rect 79 80 113 114
rect -257 -30 -223 30
rect -161 -30 -127 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 127 -30 161 30
rect 223 -30 257 30
rect -209 -114 -175 -80
rect -17 -114 17 -80
rect 175 -114 209 -80
<< metal1 >>
rect -125 114 -67 120
rect -125 80 -113 114
rect -79 80 -67 114
rect -125 74 -67 80
rect 67 114 125 120
rect 67 80 79 114
rect 113 80 125 114
rect 67 74 125 80
rect -263 30 -217 42
rect -263 -30 -257 30
rect -223 -30 -217 30
rect -263 -42 -217 -30
rect -167 30 -121 42
rect -167 -30 -161 30
rect -127 -30 -121 30
rect -167 -42 -121 -30
rect -71 30 -25 42
rect -71 -30 -65 30
rect -31 -30 -25 30
rect -71 -42 -25 -30
rect 25 30 71 42
rect 25 -30 31 30
rect 65 -30 71 30
rect 25 -42 71 -30
rect 121 30 167 42
rect 121 -30 127 30
rect 161 -30 167 30
rect 121 -42 167 -30
rect 217 30 263 42
rect 217 -30 223 30
rect 257 -30 263 30
rect 217 -42 263 -30
rect -221 -80 -163 -74
rect -221 -114 -209 -80
rect -175 -114 -163 -80
rect -221 -120 -163 -114
rect -29 -80 29 -74
rect -29 -114 -17 -80
rect 17 -114 29 -80
rect -29 -120 29 -114
rect 163 -80 221 -74
rect 163 -114 175 -80
rect 209 -114 221 -80
rect 163 -120 221 -114
<< properties >>
string FIXED_BBOX -354 -199 354 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
