magic
tech sky130A
magscale 1 2
timestamp 1717366634
<< pwell >>
rect -989 -300 989 300
<< nnmos >>
rect -761 -42 -661 42
rect -603 -42 -503 42
rect -445 -42 -345 42
rect -287 -42 -187 42
rect -129 -42 -29 42
rect 29 -42 129 42
rect 187 -42 287 42
rect 345 -42 445 42
rect 503 -42 603 42
rect 661 -42 761 42
<< mvndiff >>
rect -819 30 -761 42
rect -819 -30 -807 30
rect -773 -30 -761 30
rect -819 -42 -761 -30
rect -661 30 -603 42
rect -661 -30 -649 30
rect -615 -30 -603 30
rect -661 -42 -603 -30
rect -503 30 -445 42
rect -503 -30 -491 30
rect -457 -30 -445 30
rect -503 -42 -445 -30
rect -345 30 -287 42
rect -345 -30 -333 30
rect -299 -30 -287 30
rect -345 -42 -287 -30
rect -187 30 -129 42
rect -187 -30 -175 30
rect -141 -30 -129 30
rect -187 -42 -129 -30
rect -29 30 29 42
rect -29 -30 -17 30
rect 17 -30 29 30
rect -29 -42 29 -30
rect 129 30 187 42
rect 129 -30 141 30
rect 175 -30 187 30
rect 129 -42 187 -30
rect 287 30 345 42
rect 287 -30 299 30
rect 333 -30 345 30
rect 287 -42 345 -30
rect 445 30 503 42
rect 445 -30 457 30
rect 491 -30 503 30
rect 445 -42 503 -30
rect 603 30 661 42
rect 603 -30 615 30
rect 649 -30 661 30
rect 603 -42 661 -30
rect 761 30 819 42
rect 761 -30 773 30
rect 807 -30 819 30
rect 761 -42 819 -30
<< mvndiffc >>
rect -807 -30 -773 30
rect -649 -30 -615 30
rect -491 -30 -457 30
rect -333 -30 -299 30
rect -175 -30 -141 30
rect -17 -30 17 30
rect 141 -30 175 30
rect 299 -30 333 30
rect 457 -30 491 30
rect 615 -30 649 30
rect 773 -30 807 30
<< mvpsubdiff >>
rect -953 252 953 264
rect -953 218 -845 252
rect 845 218 953 252
rect -953 206 953 218
rect -953 156 -895 206
rect -953 -156 -941 156
rect -907 -156 -895 156
rect 895 156 953 206
rect -953 -206 -895 -156
rect 895 -156 907 156
rect 941 -156 953 156
rect 895 -206 953 -156
rect -953 -218 953 -206
rect -953 -252 -845 -218
rect 845 -252 953 -218
rect -953 -264 953 -252
<< mvpsubdiffcont >>
rect -845 218 845 252
rect -941 -156 -907 156
rect 907 -156 941 156
rect -845 -252 845 -218
<< poly >>
rect -761 114 -661 130
rect -761 80 -745 114
rect -677 80 -661 114
rect -761 42 -661 80
rect -603 114 -503 130
rect -603 80 -587 114
rect -519 80 -503 114
rect -603 42 -503 80
rect -445 114 -345 130
rect -445 80 -429 114
rect -361 80 -345 114
rect -445 42 -345 80
rect -287 114 -187 130
rect -287 80 -271 114
rect -203 80 -187 114
rect -287 42 -187 80
rect -129 114 -29 130
rect -129 80 -113 114
rect -45 80 -29 114
rect -129 42 -29 80
rect 29 114 129 130
rect 29 80 45 114
rect 113 80 129 114
rect 29 42 129 80
rect 187 114 287 130
rect 187 80 203 114
rect 271 80 287 114
rect 187 42 287 80
rect 345 114 445 130
rect 345 80 361 114
rect 429 80 445 114
rect 345 42 445 80
rect 503 114 603 130
rect 503 80 519 114
rect 587 80 603 114
rect 503 42 603 80
rect 661 114 761 130
rect 661 80 677 114
rect 745 80 761 114
rect 661 42 761 80
rect -761 -80 -661 -42
rect -761 -114 -745 -80
rect -677 -114 -661 -80
rect -761 -130 -661 -114
rect -603 -80 -503 -42
rect -603 -114 -587 -80
rect -519 -114 -503 -80
rect -603 -130 -503 -114
rect -445 -80 -345 -42
rect -445 -114 -429 -80
rect -361 -114 -345 -80
rect -445 -130 -345 -114
rect -287 -80 -187 -42
rect -287 -114 -271 -80
rect -203 -114 -187 -80
rect -287 -130 -187 -114
rect -129 -80 -29 -42
rect -129 -114 -113 -80
rect -45 -114 -29 -80
rect -129 -130 -29 -114
rect 29 -80 129 -42
rect 29 -114 45 -80
rect 113 -114 129 -80
rect 29 -130 129 -114
rect 187 -80 287 -42
rect 187 -114 203 -80
rect 271 -114 287 -80
rect 187 -130 287 -114
rect 345 -80 445 -42
rect 345 -114 361 -80
rect 429 -114 445 -80
rect 345 -130 445 -114
rect 503 -80 603 -42
rect 503 -114 519 -80
rect 587 -114 603 -80
rect 503 -130 603 -114
rect 661 -80 761 -42
rect 661 -114 677 -80
rect 745 -114 761 -80
rect 661 -130 761 -114
<< polycont >>
rect -745 80 -677 114
rect -587 80 -519 114
rect -429 80 -361 114
rect -271 80 -203 114
rect -113 80 -45 114
rect 45 80 113 114
rect 203 80 271 114
rect 361 80 429 114
rect 519 80 587 114
rect 677 80 745 114
rect -745 -114 -677 -80
rect -587 -114 -519 -80
rect -429 -114 -361 -80
rect -271 -114 -203 -80
rect -113 -114 -45 -80
rect 45 -114 113 -80
rect 203 -114 271 -80
rect 361 -114 429 -80
rect 519 -114 587 -80
rect 677 -114 745 -80
<< locali >>
rect -941 218 -845 252
rect 845 218 941 252
rect -941 156 -907 218
rect 907 156 941 218
rect -761 80 -745 114
rect -677 80 -661 114
rect -603 80 -587 114
rect -519 80 -503 114
rect -445 80 -429 114
rect -361 80 -345 114
rect -287 80 -271 114
rect -203 80 -187 114
rect -129 80 -113 114
rect -45 80 -29 114
rect 29 80 45 114
rect 113 80 129 114
rect 187 80 203 114
rect 271 80 287 114
rect 345 80 361 114
rect 429 80 445 114
rect 503 80 519 114
rect 587 80 603 114
rect 661 80 677 114
rect 745 80 761 114
rect -807 30 -773 46
rect -807 -46 -773 -30
rect -649 30 -615 46
rect -649 -46 -615 -30
rect -491 30 -457 46
rect -491 -46 -457 -30
rect -333 30 -299 46
rect -333 -46 -299 -30
rect -175 30 -141 46
rect -175 -46 -141 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 141 30 175 46
rect 141 -46 175 -30
rect 299 30 333 46
rect 299 -46 333 -30
rect 457 30 491 46
rect 457 -46 491 -30
rect 615 30 649 46
rect 615 -46 649 -30
rect 773 30 807 46
rect 773 -46 807 -30
rect -761 -114 -745 -80
rect -677 -114 -661 -80
rect -603 -114 -587 -80
rect -519 -114 -503 -80
rect -445 -114 -429 -80
rect -361 -114 -345 -80
rect -287 -114 -271 -80
rect -203 -114 -187 -80
rect -129 -114 -113 -80
rect -45 -114 -29 -80
rect 29 -114 45 -80
rect 113 -114 129 -80
rect 187 -114 203 -80
rect 271 -114 287 -80
rect 345 -114 361 -80
rect 429 -114 445 -80
rect 503 -114 519 -80
rect 587 -114 603 -80
rect 661 -114 677 -80
rect 745 -114 761 -80
rect -941 -218 -907 -156
rect 907 -218 941 -156
rect -941 -252 -845 -218
rect 845 -252 941 -218
<< viali >>
rect -745 80 -677 114
rect -587 80 -519 114
rect -429 80 -361 114
rect -271 80 -203 114
rect -113 80 -45 114
rect 45 80 113 114
rect 203 80 271 114
rect 361 80 429 114
rect 519 80 587 114
rect 677 80 745 114
rect -807 -30 -773 30
rect -649 -30 -615 30
rect -491 -30 -457 30
rect -333 -30 -299 30
rect -175 -30 -141 30
rect -17 -30 17 30
rect 141 -30 175 30
rect 299 -30 333 30
rect 457 -30 491 30
rect 615 -30 649 30
rect 773 -30 807 30
rect -745 -114 -677 -80
rect -587 -114 -519 -80
rect -429 -114 -361 -80
rect -271 -114 -203 -80
rect -113 -114 -45 -80
rect 45 -114 113 -80
rect 203 -114 271 -80
rect 361 -114 429 -80
rect 519 -114 587 -80
rect 677 -114 745 -80
<< metal1 >>
rect -757 114 -665 120
rect -757 80 -745 114
rect -677 80 -665 114
rect -757 74 -665 80
rect -599 114 -507 120
rect -599 80 -587 114
rect -519 80 -507 114
rect -599 74 -507 80
rect -441 114 -349 120
rect -441 80 -429 114
rect -361 80 -349 114
rect -441 74 -349 80
rect -283 114 -191 120
rect -283 80 -271 114
rect -203 80 -191 114
rect -283 74 -191 80
rect -125 114 -33 120
rect -125 80 -113 114
rect -45 80 -33 114
rect -125 74 -33 80
rect 33 114 125 120
rect 33 80 45 114
rect 113 80 125 114
rect 33 74 125 80
rect 191 114 283 120
rect 191 80 203 114
rect 271 80 283 114
rect 191 74 283 80
rect 349 114 441 120
rect 349 80 361 114
rect 429 80 441 114
rect 349 74 441 80
rect 507 114 599 120
rect 507 80 519 114
rect 587 80 599 114
rect 507 74 599 80
rect 665 114 757 120
rect 665 80 677 114
rect 745 80 757 114
rect 665 74 757 80
rect -813 30 -767 42
rect -813 -30 -807 30
rect -773 -30 -767 30
rect -813 -42 -767 -30
rect -655 30 -609 42
rect -655 -30 -649 30
rect -615 -30 -609 30
rect -655 -42 -609 -30
rect -497 30 -451 42
rect -497 -30 -491 30
rect -457 -30 -451 30
rect -497 -42 -451 -30
rect -339 30 -293 42
rect -339 -30 -333 30
rect -299 -30 -293 30
rect -339 -42 -293 -30
rect -181 30 -135 42
rect -181 -30 -175 30
rect -141 -30 -135 30
rect -181 -42 -135 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 135 30 181 42
rect 135 -30 141 30
rect 175 -30 181 30
rect 135 -42 181 -30
rect 293 30 339 42
rect 293 -30 299 30
rect 333 -30 339 30
rect 293 -42 339 -30
rect 451 30 497 42
rect 451 -30 457 30
rect 491 -30 497 30
rect 451 -42 497 -30
rect 609 30 655 42
rect 609 -30 615 30
rect 649 -30 655 30
rect 609 -42 655 -30
rect 767 30 813 42
rect 767 -30 773 30
rect 807 -30 813 30
rect 767 -42 813 -30
rect -757 -80 -665 -74
rect -757 -114 -745 -80
rect -677 -114 -665 -80
rect -757 -120 -665 -114
rect -599 -80 -507 -74
rect -599 -114 -587 -80
rect -519 -114 -507 -80
rect -599 -120 -507 -114
rect -441 -80 -349 -74
rect -441 -114 -429 -80
rect -361 -114 -349 -80
rect -441 -120 -349 -114
rect -283 -80 -191 -74
rect -283 -114 -271 -80
rect -203 -114 -191 -80
rect -283 -120 -191 -114
rect -125 -80 -33 -74
rect -125 -114 -113 -80
rect -45 -114 -33 -80
rect -125 -120 -33 -114
rect 33 -80 125 -74
rect 33 -114 45 -80
rect 113 -114 125 -80
rect 33 -120 125 -114
rect 191 -80 283 -74
rect 191 -114 203 -80
rect 271 -114 283 -80
rect 191 -120 283 -114
rect 349 -80 441 -74
rect 349 -114 361 -80
rect 429 -114 441 -80
rect 349 -120 441 -114
rect 507 -80 599 -74
rect 507 -114 519 -80
rect 587 -114 599 -80
rect 507 -120 599 -114
rect 665 -80 757 -74
rect 665 -114 677 -80
rect 745 -114 757 -80
rect 665 -120 757 -114
<< properties >>
string FIXED_BBOX -924 -235 924 235
string gencell sky130_fd_pr__nfet_03v3_nvt
string library sky130
string parameters w 0.42 l 0.5 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
