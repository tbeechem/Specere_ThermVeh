magic
tech sky130A
magscale 1 2
timestamp 1717349526
<< pwell >>
rect 32 -514 986 -265
rect 1000 -492 1070 -374
rect 1282 -490 1352 -372
rect 32 -792 572 -514
rect 608 -792 986 -514
rect 998 -716 1094 -644
rect 1288 -706 1352 -652
rect 1514 -684 1546 -520
rect 1288 -716 1350 -706
rect 996 -758 1350 -716
rect 32 -865 986 -792
<< locali >>
rect -16 -384 1352 -348
rect -16 -720 20 -384
rect 184 -490 254 -384
rect 452 -490 522 -384
rect 1000 -492 1070 -384
rect 1282 -490 1352 -384
rect 442 -720 536 -646
rect 998 -716 1094 -644
rect 1288 -706 1352 -652
rect 1288 -716 1350 -706
rect 996 -720 1350 -716
rect -16 -722 1350 -720
rect -16 -756 200 -722
rect 238 -756 1350 -722
rect 996 -758 1350 -756
<< viali >>
rect 200 -756 238 -722
<< metal1 >>
rect 0 -150 200 50
rect 672 -122 850 50
rect 98 -356 128 -150
rect 672 -182 718 -122
rect 812 -182 850 -122
rect 1350 -150 1550 50
rect 672 -216 850 -182
rect 98 -384 1248 -356
rect 98 -598 128 -384
rect 292 -554 326 -520
rect 178 -680 182 -644
rect 178 -722 246 -680
rect 178 -756 200 -722
rect 238 -756 246 -722
rect 178 -900 246 -756
rect 292 -791 328 -554
rect 378 -791 414 -518
rect 570 -626 604 -384
rect 648 -628 682 -384
rect 714 -424 816 -416
rect 714 -482 722 -424
rect 808 -482 816 -424
rect 714 -490 816 -482
rect 714 -648 816 -640
rect 714 -706 722 -648
rect 808 -706 816 -648
rect 714 -714 816 -706
rect 292 -792 572 -791
rect 850 -792 888 -522
rect 924 -792 962 -524
rect 1128 -626 1162 -384
rect 1198 -622 1232 -384
rect 1514 -522 1548 -150
rect 1394 -532 1548 -522
rect 1394 -592 1546 -532
rect 1514 -644 1546 -592
rect 1514 -792 1550 -644
rect 292 -794 1550 -792
rect 294 -824 1550 -794
rect 294 -825 862 -824
rect 294 -828 328 -825
rect 570 -826 862 -825
rect 150 -1100 350 -900
rect 672 -976 850 -940
rect 672 -1036 716 -976
rect 810 -1036 850 -976
rect 672 -1206 850 -1036
<< via1 >>
rect 718 -182 812 -122
rect 722 -482 808 -424
rect 722 -706 808 -648
rect 716 -1036 810 -976
<< metal2 >>
rect 678 -122 850 -102
rect 678 -182 718 -122
rect 812 -182 850 -122
rect 678 -210 850 -182
rect 714 -424 816 -210
rect 714 -482 722 -424
rect 808 -482 816 -424
rect 714 -488 816 -482
rect 714 -648 816 -644
rect 714 -706 722 -648
rect 808 -706 816 -648
rect 714 -952 816 -706
rect 674 -976 846 -952
rect 674 -1036 716 -976
rect 810 -1036 846 -976
rect 674 -1060 846 -1036
use sky130_fd_pr__nfet_03v3_nvt_VB5P9F  sky130_fd_pr__nfet_03v3_nvt_VB5P9F_0
timestamp 1717306961
transform 1 0 765 0 1 -565
box -830 -300 830 300
<< labels >>
flabel metal1 0 -150 200 50 0 FreeSans 256 0 0 0 VD_H
port 0 nsew
flabel metal1 150 -1100 350 -900 0 FreeSans 256 0 0 0 VG_H
port 1 nsew
flabel metal1 1350 -150 1550 50 0 FreeSans 256 0 0 0 VLow_Src
port 2 nsew
<< end >>
