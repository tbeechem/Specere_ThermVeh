magic
tech sky130A
timestamp 1717306961
<< pwell >>
rect -297 -150 297 150
<< nnmos >>
rect -183 -21 -133 21
rect -104 -21 -54 21
rect -25 -21 25 21
rect 54 -21 104 21
rect 133 -21 183 21
<< mvndiff >>
rect -212 15 -183 21
rect -212 -15 -206 15
rect -189 -15 -183 15
rect -212 -21 -183 -15
rect -133 15 -104 21
rect -133 -15 -127 15
rect -110 -15 -104 15
rect -133 -21 -104 -15
rect -54 15 -25 21
rect -54 -15 -48 15
rect -31 -15 -25 15
rect -54 -21 -25 -15
rect 25 15 54 21
rect 25 -15 31 15
rect 48 -15 54 15
rect 25 -21 54 -15
rect 104 15 133 21
rect 104 -15 110 15
rect 127 -15 133 15
rect 104 -21 133 -15
rect 183 15 212 21
rect 183 -15 189 15
rect 206 -15 212 15
rect 183 -21 212 -15
<< mvndiffc >>
rect -206 -15 -189 15
rect -127 -15 -110 15
rect -48 -15 -31 15
rect 31 -15 48 15
rect 110 -15 127 15
rect 189 -15 206 15
<< mvpsubdiff >>
rect -279 126 279 132
rect -279 109 -225 126
rect 225 109 279 126
rect -279 103 279 109
rect -279 78 -250 103
rect -279 -78 -273 78
rect -256 -78 -250 78
rect 250 78 279 103
rect -279 -103 -250 -78
rect 250 -78 256 78
rect 273 -78 279 78
rect 250 -103 279 -78
rect -279 -109 279 -103
rect -279 -126 -225 -109
rect 225 -126 279 -109
rect -279 -132 279 -126
<< mvpsubdiffcont >>
rect -225 109 225 126
rect -273 -78 -256 78
rect 256 -78 273 78
rect -225 -126 225 -109
<< poly >>
rect -183 57 -133 65
rect -183 40 -175 57
rect -141 40 -133 57
rect -183 21 -133 40
rect -104 57 -54 65
rect -104 40 -96 57
rect -62 40 -54 57
rect -104 21 -54 40
rect -25 57 25 65
rect -25 40 -17 57
rect 17 40 25 57
rect -25 21 25 40
rect 54 57 104 65
rect 54 40 62 57
rect 96 40 104 57
rect 54 21 104 40
rect 133 57 183 65
rect 133 40 141 57
rect 175 40 183 57
rect 133 21 183 40
rect -183 -40 -133 -21
rect -183 -57 -175 -40
rect -141 -57 -133 -40
rect -183 -65 -133 -57
rect -104 -40 -54 -21
rect -104 -57 -96 -40
rect -62 -57 -54 -40
rect -104 -65 -54 -57
rect -25 -40 25 -21
rect -25 -57 -17 -40
rect 17 -57 25 -40
rect -25 -65 25 -57
rect 54 -40 104 -21
rect 54 -57 62 -40
rect 96 -57 104 -40
rect 54 -65 104 -57
rect 133 -40 183 -21
rect 133 -57 141 -40
rect 175 -57 183 -40
rect 133 -65 183 -57
<< polycont >>
rect -175 40 -141 57
rect -96 40 -62 57
rect -17 40 17 57
rect 62 40 96 57
rect 141 40 175 57
rect -175 -57 -141 -40
rect -96 -57 -62 -40
rect -17 -57 17 -40
rect 62 -57 96 -40
rect 141 -57 175 -40
<< locali >>
rect -273 109 -225 126
rect 225 109 273 126
rect -273 78 -256 109
rect 256 78 273 109
rect -183 40 -175 57
rect -141 40 -133 57
rect -104 40 -96 57
rect -62 40 -54 57
rect -25 40 -17 57
rect 17 40 25 57
rect 54 40 62 57
rect 96 40 104 57
rect 133 40 141 57
rect 175 40 183 57
rect -206 15 -189 23
rect -206 -23 -189 -15
rect -127 15 -110 23
rect -127 -23 -110 -15
rect -48 15 -31 23
rect -48 -23 -31 -15
rect 31 15 48 23
rect 31 -23 48 -15
rect 110 15 127 23
rect 110 -23 127 -15
rect 189 15 206 23
rect 189 -23 206 -15
rect -183 -57 -175 -40
rect -141 -57 -133 -40
rect -104 -57 -96 -40
rect -62 -57 -54 -40
rect -25 -57 -17 -40
rect 17 -57 25 -40
rect 54 -57 62 -40
rect 96 -57 104 -40
rect 133 -57 141 -40
rect 175 -57 183 -40
rect -273 -109 -256 -78
rect 256 -109 273 -78
rect -273 -126 -225 -109
rect 225 -126 273 -109
<< viali >>
rect -175 40 -141 57
rect -96 40 -62 57
rect -17 40 17 57
rect 62 40 96 57
rect 141 40 175 57
rect -206 -15 -189 15
rect -127 -15 -110 15
rect -48 -15 -31 15
rect 31 -15 48 15
rect 110 -15 127 15
rect 189 -15 206 15
rect -175 -57 -141 -40
rect -96 -57 -62 -40
rect -17 -57 17 -40
rect 62 -57 96 -40
rect 141 -57 175 -40
<< metal1 >>
rect -181 57 -135 60
rect -181 40 -175 57
rect -141 40 -135 57
rect -181 37 -135 40
rect -102 57 -56 60
rect -102 40 -96 57
rect -62 40 -56 57
rect -102 37 -56 40
rect -23 57 23 60
rect -23 40 -17 57
rect 17 40 23 57
rect -23 37 23 40
rect 56 57 102 60
rect 56 40 62 57
rect 96 40 102 57
rect 56 37 102 40
rect 135 57 181 60
rect 135 40 141 57
rect 175 40 181 57
rect 135 37 181 40
rect -209 15 -186 21
rect -209 -15 -206 15
rect -189 -15 -186 15
rect -209 -21 -186 -15
rect -130 15 -107 21
rect -130 -15 -127 15
rect -110 -15 -107 15
rect -130 -21 -107 -15
rect -51 15 -28 21
rect -51 -15 -48 15
rect -31 -15 -28 15
rect -51 -21 -28 -15
rect 28 15 51 21
rect 28 -15 31 15
rect 48 -15 51 15
rect 28 -21 51 -15
rect 107 15 130 21
rect 107 -15 110 15
rect 127 -15 130 15
rect 107 -21 130 -15
rect 186 15 209 21
rect 186 -15 189 15
rect 206 -15 209 15
rect 186 -21 209 -15
rect -181 -40 -135 -37
rect -181 -57 -175 -40
rect -141 -57 -135 -40
rect -181 -60 -135 -57
rect -102 -40 -56 -37
rect -102 -57 -96 -40
rect -62 -57 -56 -40
rect -102 -60 -56 -57
rect -23 -40 23 -37
rect -23 -57 -17 -40
rect 17 -57 23 -40
rect -23 -60 23 -57
rect 56 -40 102 -37
rect 56 -57 62 -40
rect 96 -57 102 -40
rect 56 -60 102 -57
rect 135 -40 181 -37
rect 135 -57 141 -40
rect 175 -57 181 -40
rect 135 -60 181 -57
<< properties >>
string FIXED_BBOX -264 -117 264 117
string gencell sky130_fd_pr__nfet_03v3_nvt
string library sky130
string parameters w 0.42 l 0.5 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
