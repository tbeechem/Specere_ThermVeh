magic
tech sky130A
magscale 1 2
timestamp 1717296424
<< metal1 >>
rect -800 -450 -600 -400
rect 900 -450 1100 -400
rect -800 -550 150 -450
rect 300 -550 1100 -450
rect -800 -600 -600 -550
rect 900 -600 1100 -550
rect 150 -1100 250 -650
rect 100 -1300 300 -1100
use sky130_fd_pr__nfet_03v3_nvt_EJ4KLV  XM1
timestamp 1717296329
transform 1 0 213 0 1 -507
box -278 -358 278 358
<< labels >>
flabel metal1 -800 -600 -600 -400 0 FreeSans 160 0 0 0 VD_H
port 0 nsew
flabel metal1 900 -600 1100 -400 0 FreeSans 160 0 0 0 VLow_Src
port 2 nsew
flabel metal1 100 -1300 300 -1100 0 FreeSans 160 0 0 0 VG_H
port 1 nsew
<< end >>
