magic
tech sky130A
magscale 1 2
timestamp 1717386517
<< metal1 >>
rect 5996 12654 7448 13018
rect 5996 11830 6392 12654
rect 7118 11830 7448 12654
rect 5996 2973 7448 11830
rect -7965 650 -7017 656
rect -7965 -1342 -7017 -298
rect 9210 -1068 10694 -983
rect 9193 -2006 10694 -1068
rect -5363 -2521 -1549 -2321
rect -5363 -4752 -5163 -2521
rect 9193 -3513 10694 -3507
rect -6088 -11910 -4636 -4752
rect -6088 -12734 -5758 -11910
rect -5032 -12734 -4636 -11910
rect -6088 -13328 -4636 -12734
<< via1 >>
rect 6392 11830 7118 12654
rect -7965 -298 -7017 650
rect 9193 -3507 10694 -2006
rect -5758 -12734 -5032 -11910
<< metal2 >>
rect 6030 14670 7350 15100
rect 6030 13944 6392 14670
rect 7084 13944 7350 14670
rect 6030 12654 7350 13944
rect 6030 11830 6392 12654
rect 7118 11830 7350 12654
rect 6030 11468 7350 11830
rect -1260 6240 -300 6360
rect -1260 5580 -1080 6240
rect -420 5580 -300 6240
rect -1260 3703 -300 5580
rect 2460 6240 3420 6360
rect 2460 5580 2640 6240
rect 3300 5580 3420 6240
rect 2460 3703 3420 5580
rect -2615 3142 3421 3703
rect -7974 1355 -7965 2303
rect -7017 1355 -7008 2303
rect -7965 650 -7017 1355
rect -7971 -298 -7965 650
rect -7017 -298 -7011 650
rect -2615 -372 -2054 3142
rect -1260 3138 -300 3142
rect 2460 3121 3420 3142
rect -2937 -3623 -2598 -2273
rect 9187 -3507 9193 -2006
rect 10694 -3507 10700 -2006
rect -1320 -3623 -360 -3615
rect 2400 -3623 3345 -3593
rect -2937 -3962 3345 -3623
rect -2937 -3988 -2598 -3962
rect -1320 -6240 -360 -3962
rect -1320 -6900 -1140 -6240
rect -480 -6900 -360 -6240
rect -1320 -7020 -360 -6900
rect 2400 -4328 3345 -3962
rect 9193 -4052 10694 -3507
rect 2400 -6240 3360 -4328
rect 9193 -5562 10694 -5553
rect 2400 -6900 2580 -6240
rect 3240 -6900 3360 -6240
rect 2400 -7020 3360 -6900
rect -6054 -11910 -4734 -11742
rect -6054 -12734 -5758 -11910
rect -5032 -12734 -4734 -11910
rect -6054 -14352 -4734 -12734
rect -6054 -15078 -5790 -14352
rect -5098 -15078 -4734 -14352
rect -6054 -15374 -4734 -15078
<< via2 >>
rect 6392 13944 7084 14670
rect -1080 5580 -420 6240
rect 2640 5580 3300 6240
rect -7965 1355 -7017 2303
rect -1140 -6900 -480 -6240
rect 9193 -5553 10694 -4052
rect 2580 -6900 3240 -6240
rect -5790 -15078 -5098 -14352
<< metal3 >>
rect 6126 17284 7316 17692
rect 6126 16360 6352 17284
rect 7028 16360 7316 17284
rect 6126 14670 7316 16360
rect 6126 13944 6392 14670
rect 7084 13944 7316 14670
rect 6126 13596 7316 13944
rect -1260 9240 -300 9480
rect -1260 8460 -1080 9240
rect -420 8460 -300 9240
rect -1260 6240 -300 8460
rect -1260 5580 -1080 6240
rect -420 5580 -300 6240
rect -1260 5400 -300 5580
rect 2460 9240 3420 9480
rect 2460 8460 2640 9240
rect 3300 8460 3420 9240
rect 2460 6240 3420 8460
rect 2460 5580 2640 6240
rect 3300 5580 3420 6240
rect 2460 5400 3420 5580
rect -7970 2303 -7012 2308
rect -9353 1355 -9347 2303
rect -8399 1355 -7965 2303
rect -7017 1355 -7012 2303
rect -7970 1350 -7012 1355
rect 9188 -4051 10699 -4047
rect 9188 -4052 11427 -4051
rect 9188 -5553 9193 -4052
rect 10694 -5552 11427 -4052
rect 12928 -5552 12934 -4051
rect 10694 -5553 10699 -5552
rect 9188 -5558 10699 -5553
rect -1320 -6240 -360 -6060
rect -1320 -6900 -1140 -6240
rect -480 -6900 -360 -6240
rect -1320 -9120 -360 -6900
rect -1320 -9900 -1140 -9120
rect -480 -9900 -360 -9120
rect -1320 -10140 -360 -9900
rect 2400 -6240 3360 -6060
rect 2400 -6900 2580 -6240
rect 3240 -6900 3360 -6240
rect 2400 -9120 3360 -6900
rect 2400 -9900 2580 -9120
rect 3240 -9900 3360 -9120
rect 2400 -10140 3360 -9900
rect -6054 -14352 -4864 -14150
rect -6054 -15078 -5790 -14352
rect -5098 -15078 -4864 -14352
rect -6054 -17042 -4864 -15078
rect -6054 -17966 -5794 -17042
rect -5118 -17966 -4864 -17042
rect -6054 -18246 -4864 -17966
<< via3 >>
rect 6352 16360 7028 17284
rect -1080 8460 -420 9240
rect 2640 8460 3300 9240
rect -9347 1355 -8399 2303
rect 11427 -5552 12928 -4051
rect -1140 -9900 -480 -9120
rect 2580 -9900 3240 -9120
rect -5794 -17966 -5118 -17042
<< metal4 >>
rect 5418 24654 7998 25298
rect 5418 22976 5934 24654
rect 7354 22976 7998 24654
rect 5418 17284 7998 22976
rect 5418 16360 6352 17284
rect 7028 16360 7998 17284
rect 5418 15752 7998 16360
rect -1260 12660 -300 12900
rect -1260 12180 -1140 12660
rect -420 12180 -300 12660
rect -1260 9240 -300 12180
rect -1260 8460 -1080 9240
rect -420 8460 -300 9240
rect -1260 8100 -300 8460
rect 2460 12660 3420 12900
rect 2460 12180 2580 12660
rect 3300 12180 3420 12660
rect 2460 9240 3420 12180
rect 2460 8460 2640 9240
rect 3300 8460 3420 9240
rect 2460 8100 3420 8460
rect -9348 2303 -8398 2304
rect -10729 1355 -9347 2303
rect -8399 1355 -8398 2303
rect -10729 -366 -9781 1355
rect -9348 1354 -8398 1355
rect 11427 -4050 12928 -1478
rect 11426 -4051 12929 -4050
rect 11426 -5552 11427 -4051
rect 12928 -5552 12929 -4051
rect 11426 -5553 12929 -5552
rect -1320 -9120 -360 -8760
rect -1320 -9900 -1140 -9120
rect -480 -9900 -360 -9120
rect -1320 -12840 -360 -9900
rect -1320 -13320 -1200 -12840
rect -480 -13320 -360 -12840
rect -1320 -13560 -360 -13320
rect 2400 -9120 3360 -8760
rect 2400 -9900 2580 -9120
rect 3240 -9900 3360 -9120
rect 2400 -12840 3360 -9900
rect 2400 -13320 2520 -12840
rect 3240 -13320 3360 -12840
rect 2400 -13560 3360 -13320
rect -6644 -17042 -4064 -16694
rect -6644 -17966 -5794 -17042
rect -5118 -17966 -4064 -17042
rect -6644 -23918 -4064 -17966
rect -6644 -25596 -6064 -23918
rect -4644 -25596 -4064 -23918
rect -6644 -26240 -4064 -25596
<< via4 >>
rect 5934 22976 7354 24654
rect -1140 12180 -420 12660
rect 2580 12180 3300 12660
rect -10729 -1314 -9781 -366
rect 11427 -1478 12928 23
rect -1200 -13320 -480 -12840
rect 2520 -13320 3240 -12840
rect -6064 -25596 -4644 -23918
<< metal5 >>
rect -7104 25824 8896 42024
rect -28066 20160 -12066 25780
rect 5418 24654 7978 25824
rect 5418 22976 5934 24654
rect 7354 22976 7978 24654
rect 5418 22068 7978 22976
rect -28066 18900 -300 20160
rect 15120 20100 31120 25800
rect 14160 20084 31120 20100
rect 2392 18968 31120 20084
rect 2392 18952 5438 18968
rect 14160 18960 31120 18968
rect -28066 17000 -12066 18900
rect -28200 16000 -12060 17000
rect -28066 9580 -12066 16000
rect -1274 13080 -306 18900
rect -1294 12660 -284 13080
rect -1294 12180 -1140 12660
rect -420 12180 -284 12660
rect -1294 11980 -284 12180
rect 2426 12660 3436 18952
rect 2426 12180 2580 12660
rect 3300 12180 3436 12660
rect 2426 11980 3436 12180
rect 15120 9600 31120 18960
rect -28000 -86 -12000 7100
rect 15030 54 31030 7066
rect 11403 24 12952 47
rect 14351 24 31030 54
rect 11403 23 31030 24
rect -28000 -361 -11982 -86
rect -28000 -366 -11624 -361
rect -10753 -366 -9757 -342
rect -28000 -1314 -10729 -366
rect -9781 -1314 -9757 -366
rect -28000 -1315 -11624 -1314
rect -28000 -1376 -11996 -1315
rect -10753 -1338 -9757 -1314
rect -28000 -9100 -12000 -1376
rect 11403 -1478 11427 23
rect 12928 -1477 31030 23
rect 12928 -1478 12952 -1477
rect 11403 -1502 12952 -1478
rect 14351 -1486 31030 -1477
rect 15030 -9134 31030 -1486
rect -28080 -19776 -12080 -11622
rect -1354 -12840 -344 -12640
rect -1354 -13320 -1200 -12840
rect -480 -13320 -344 -12840
rect -1354 -13740 -344 -13320
rect 2366 -12840 3376 -12640
rect 2366 -13320 2520 -12840
rect 3240 -13320 3376 -12840
rect -1334 -19776 -366 -13740
rect 2366 -19612 3376 -13320
rect 2332 -19628 5378 -19612
rect 15030 -19628 31030 -11764
rect -28080 -20702 -326 -19776
rect -28080 -27822 -12080 -20702
rect 2332 -20744 31030 -19628
rect 15002 -20852 31030 -20744
rect -6592 -23918 -4032 -23134
rect -6592 -25596 -6064 -23918
rect -4644 -25596 -4032 -23918
rect -6592 -27864 -4032 -25596
rect -7616 -44064 8384 -27864
rect 15030 -27964 31030 -20852
<< glass >>
rect -6800 26200 8600 41600
rect -27600 9800 -12466 25380
rect 15520 10000 30600 25400
rect -27600 -8700 -12400 6700
rect 15430 -8734 30630 6666
rect -27680 -27400 -12480 -12020
rect 15430 -27564 30630 -12164
rect -7200 -43800 8000 -28200
use GSense_nFET_6Contacts_V2  GSense_nFET_3VD_3Vg_5nf_V2_0 ~/Specere_ThermVeh/mag
timestamp 1717352107
transform 1 0 315 0 1 -138
box 0 0 1 1
use GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline  GSense_nFET_3VD_3Vg_51nf_V2AllGates_Mid_Therm_0
timestamp 1717386517
transform 1 0 -5867 0 1 -731
box -1366 -1870 15678 395
<< end >>
