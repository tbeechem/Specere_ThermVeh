magic
tech sky130A
magscale 1 2
timestamp 1717259173
<< error_p >>
rect -221 353 -220 397
rect -193 379 -192 419
<< nwell >>
rect -338 -497 338 497
<< mvpmos >>
rect -80 -200 80 200
<< mvpdiff >>
rect -138 187 -80 200
rect -138 153 -126 187
rect -92 153 -80 187
rect -138 119 -80 153
rect -138 85 -126 119
rect -92 85 -80 119
rect -138 51 -80 85
rect -138 17 -126 51
rect -92 17 -80 51
rect -138 -17 -80 17
rect -138 -51 -126 -17
rect -92 -51 -80 -17
rect -138 -85 -80 -51
rect -138 -119 -126 -85
rect -92 -119 -80 -85
rect -138 -153 -80 -119
rect -138 -187 -126 -153
rect -92 -187 -80 -153
rect -138 -200 -80 -187
rect 80 187 138 200
rect 80 153 92 187
rect 126 153 138 187
rect 80 119 138 153
rect 80 85 92 119
rect 126 85 138 119
rect 80 51 138 85
rect 80 17 92 51
rect 126 17 138 51
rect 80 -17 138 17
rect 80 -51 92 -17
rect 126 -51 138 -17
rect 80 -85 138 -51
rect 80 -119 92 -85
rect 126 -119 138 -85
rect 80 -153 138 -119
rect 80 -187 92 -153
rect 126 -187 138 -153
rect 80 -200 138 -187
<< mvpdiffc >>
rect -126 153 -92 187
rect -126 85 -92 119
rect -126 17 -92 51
rect -126 -51 -92 -17
rect -126 -119 -92 -85
rect -126 -187 -92 -153
rect 92 153 126 187
rect 92 85 126 119
rect 92 17 126 51
rect 92 -51 126 -17
rect 92 -119 126 -85
rect 92 -187 126 -153
<< mvnsubdiff >>
rect -272 419 272 431
rect -272 385 -153 419
rect -119 385 -85 419
rect -51 385 -17 419
rect 17 385 51 419
rect 85 385 119 419
rect 153 385 272 419
rect -272 373 272 385
rect -272 323 -214 373
rect -272 289 -260 323
rect -226 289 -214 323
rect 214 323 272 373
rect -272 255 -214 289
rect -272 221 -260 255
rect -226 221 -214 255
rect -272 187 -214 221
rect 214 289 226 323
rect 260 289 272 323
rect 214 255 272 289
rect 214 221 226 255
rect 260 221 272 255
rect -272 153 -260 187
rect -226 153 -214 187
rect -272 119 -214 153
rect -272 85 -260 119
rect -226 85 -214 119
rect -272 51 -214 85
rect -272 17 -260 51
rect -226 17 -214 51
rect -272 -17 -214 17
rect -272 -51 -260 -17
rect -226 -51 -214 -17
rect -272 -85 -214 -51
rect -272 -119 -260 -85
rect -226 -119 -214 -85
rect -272 -153 -214 -119
rect -272 -187 -260 -153
rect -226 -187 -214 -153
rect -272 -221 -214 -187
rect 214 187 272 221
rect 214 153 226 187
rect 260 153 272 187
rect 214 119 272 153
rect 214 85 226 119
rect 260 85 272 119
rect 214 51 272 85
rect 214 17 226 51
rect 260 17 272 51
rect 214 -17 272 17
rect 214 -51 226 -17
rect 260 -51 272 -17
rect 214 -85 272 -51
rect 214 -119 226 -85
rect 260 -119 272 -85
rect 214 -153 272 -119
rect 214 -187 226 -153
rect 260 -187 272 -153
rect -272 -255 -260 -221
rect -226 -255 -214 -221
rect -272 -289 -214 -255
rect -272 -323 -260 -289
rect -226 -323 -214 -289
rect 214 -221 272 -187
rect 214 -255 226 -221
rect 260 -255 272 -221
rect 214 -289 272 -255
rect -272 -373 -214 -323
rect 214 -323 226 -289
rect 260 -323 272 -289
rect 214 -373 272 -323
rect -272 -385 272 -373
rect -272 -419 -153 -385
rect -119 -419 -85 -385
rect -51 -419 -17 -385
rect 17 -419 51 -385
rect 85 -419 119 -385
rect 153 -419 272 -385
rect -272 -431 272 -419
<< mvnsubdiffcont >>
rect -153 385 -119 419
rect -85 385 -51 419
rect -17 385 17 419
rect 51 385 85 419
rect 119 385 153 419
rect -260 289 -226 323
rect -260 221 -226 255
rect 226 289 260 323
rect 226 221 260 255
rect -260 153 -226 187
rect -260 85 -226 119
rect -260 17 -226 51
rect -260 -51 -226 -17
rect -260 -119 -226 -85
rect -260 -187 -226 -153
rect 226 153 260 187
rect 226 85 260 119
rect 226 17 260 51
rect 226 -51 260 -17
rect 226 -119 260 -85
rect 226 -187 260 -153
rect -260 -255 -226 -221
rect -260 -323 -226 -289
rect 226 -255 260 -221
rect 226 -323 260 -289
rect -153 -419 -119 -385
rect -85 -419 -51 -385
rect -17 -419 17 -385
rect 51 -419 85 -385
rect 119 -419 153 -385
<< poly >>
rect -80 281 80 297
rect -80 247 -51 281
rect -17 247 17 281
rect 51 247 80 281
rect -80 200 80 247
rect -80 -247 80 -200
rect -80 -281 -51 -247
rect -17 -281 17 -247
rect 51 -281 80 -247
rect -80 -297 80 -281
<< polycont >>
rect -51 247 -17 281
rect 17 247 51 281
rect -51 -281 -17 -247
rect 17 -281 51 -247
<< locali >>
rect -260 385 -161 419
rect -119 385 -89 419
rect -51 385 -17 419
rect 17 385 51 419
rect 89 385 119 419
rect 161 385 260 419
rect -260 353 -226 385
rect -260 281 -226 289
rect 226 323 260 385
rect -80 247 -53 281
rect -17 247 17 281
rect 53 247 80 281
rect 226 255 260 289
rect -260 209 -226 221
rect -260 137 -226 153
rect -260 65 -226 85
rect -260 -17 -226 17
rect -260 -85 -226 -51
rect -260 -153 -226 -119
rect -260 -221 -226 -187
rect -126 187 -92 204
rect -126 119 -92 127
rect -126 51 -92 55
rect -126 -55 -92 -51
rect -126 -127 -92 -119
rect -126 -204 -92 -187
rect 92 187 126 204
rect 92 119 126 127
rect 92 51 126 55
rect 92 -55 126 -51
rect 92 -127 126 -119
rect 92 -204 126 -187
rect 226 187 260 221
rect 226 119 260 153
rect 226 51 260 85
rect 226 -17 260 17
rect 226 -85 260 -51
rect 226 -153 260 -119
rect 226 -221 260 -187
rect -260 -289 -226 -255
rect -80 -281 -53 -247
rect -17 -281 17 -247
rect 53 -281 80 -247
rect -260 -385 -226 -323
rect 226 -289 260 -255
rect 226 -385 260 -323
rect -260 -419 -153 -385
rect -119 -419 -85 -385
rect -51 -419 -17 -385
rect 17 -419 51 -385
rect 85 -419 119 -385
rect 153 -419 260 -385
<< viali >>
rect -161 385 -153 419
rect -153 385 -127 419
rect -89 385 -85 419
rect -85 385 -55 419
rect -17 385 17 419
rect 55 385 85 419
rect 85 385 89 419
rect 127 385 153 419
rect 153 385 161 419
rect -260 323 -226 353
rect -260 319 -226 323
rect -260 255 -226 281
rect -260 247 -226 255
rect -53 247 -51 281
rect -51 247 -19 281
rect 19 247 51 281
rect 51 247 53 281
rect -260 187 -226 209
rect -260 175 -226 187
rect -260 119 -226 137
rect -260 103 -226 119
rect -260 51 -226 65
rect -260 31 -226 51
rect -126 153 -92 161
rect -126 127 -92 153
rect -126 85 -92 89
rect -126 55 -92 85
rect -126 -17 -92 17
rect -126 -85 -92 -55
rect -126 -89 -92 -85
rect -126 -153 -92 -127
rect -126 -161 -92 -153
rect 92 153 126 161
rect 92 127 126 153
rect 92 85 126 89
rect 92 55 126 85
rect 92 -17 126 17
rect 92 -85 126 -55
rect 92 -89 126 -85
rect 92 -153 126 -127
rect 92 -161 126 -153
rect -53 -281 -51 -247
rect -51 -281 -19 -247
rect 19 -281 51 -247
rect 51 -281 53 -247
<< metal1 >>
rect -193 419 193 425
rect -266 353 -220 397
rect -193 385 -161 419
rect -127 385 -89 419
rect -55 385 -17 419
rect 17 385 55 419
rect 89 385 127 419
rect 161 385 193 419
rect -193 379 193 385
rect -266 319 -260 353
rect -226 319 -220 353
rect -266 281 -220 319
rect -266 247 -260 281
rect -226 247 -220 281
rect -266 209 -220 247
rect -76 281 76 287
rect -76 247 -53 281
rect -19 247 19 281
rect 53 247 76 281
rect -76 241 76 247
rect -266 175 -260 209
rect -226 175 -220 209
rect -266 137 -220 175
rect -266 103 -260 137
rect -226 103 -220 137
rect -266 65 -220 103
rect -266 31 -260 65
rect -226 31 -220 65
rect -266 -12 -220 31
rect -132 161 -86 200
rect -132 127 -126 161
rect -92 127 -86 161
rect -132 89 -86 127
rect -132 55 -126 89
rect -92 55 -86 89
rect -132 17 -86 55
rect -132 -17 -126 17
rect -92 -17 -86 17
rect -132 -55 -86 -17
rect -132 -89 -126 -55
rect -92 -89 -86 -55
rect -132 -127 -86 -89
rect -132 -161 -126 -127
rect -92 -161 -86 -127
rect -132 -200 -86 -161
rect 86 161 132 200
rect 86 127 92 161
rect 126 127 132 161
rect 86 89 132 127
rect 86 55 92 89
rect 126 55 132 89
rect 86 17 132 55
rect 86 -17 92 17
rect 126 -17 132 17
rect 86 -55 132 -17
rect 86 -89 92 -55
rect 126 -89 132 -55
rect 86 -127 132 -89
rect 86 -161 92 -127
rect 126 -161 132 -127
rect 86 -200 132 -161
rect -76 -247 76 -241
rect -76 -281 -53 -247
rect -19 -281 19 -247
rect 53 -281 76 -247
rect -76 -287 76 -281
<< properties >>
string FIXED_BBOX -243 -402 243 402
<< end >>
