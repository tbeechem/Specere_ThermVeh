// sch_path: /home/parallels/Specere_ThermVeh/xschem/GSense_nFET_1f1WL150n_V1.sch
module GSense_nFET_1f1WL150n_V1
(
  inout wire VG_H,
  inout wire VD_H,
  inout wire VLow_Src
);
X M3  VD_H  ,  VG_H  ,  VLow_Src  ,  VLow_Src  sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
endmodule
