magic
tech sky130A
timestamp 1717306961
<< pwell >>
rect -415 -150 415 150
<< nnmos >>
rect -301 -21 -251 21
rect -163 -21 -113 21
rect -25 -21 25 21
rect 113 -21 163 21
rect 251 -21 301 21
<< mvndiff >>
rect -330 15 -301 21
rect -330 -15 -324 15
rect -307 -15 -301 15
rect -330 -21 -301 -15
rect -251 15 -222 21
rect -251 -15 -245 15
rect -228 -15 -222 15
rect -251 -21 -222 -15
rect -192 15 -163 21
rect -192 -15 -186 15
rect -169 -15 -163 15
rect -192 -21 -163 -15
rect -113 15 -84 21
rect -113 -15 -107 15
rect -90 -15 -84 15
rect -113 -21 -84 -15
rect -54 15 -25 21
rect -54 -15 -48 15
rect -31 -15 -25 15
rect -54 -21 -25 -15
rect 25 15 54 21
rect 25 -15 31 15
rect 48 -15 54 15
rect 25 -21 54 -15
rect 84 15 113 21
rect 84 -15 90 15
rect 107 -15 113 15
rect 84 -21 113 -15
rect 163 15 192 21
rect 163 -15 169 15
rect 186 -15 192 15
rect 163 -21 192 -15
rect 222 15 251 21
rect 222 -15 228 15
rect 245 -15 251 15
rect 222 -21 251 -15
rect 301 15 330 21
rect 301 -15 307 15
rect 324 -15 330 15
rect 301 -21 330 -15
<< mvndiffc >>
rect -324 -15 -307 15
rect -245 -15 -228 15
rect -186 -15 -169 15
rect -107 -15 -90 15
rect -48 -15 -31 15
rect 31 -15 48 15
rect 90 -15 107 15
rect 169 -15 186 15
rect 228 -15 245 15
rect 307 -15 324 15
<< mvpsubdiff >>
rect -397 103 397 132
rect -397 -103 -368 103
rect 368 78 397 103
rect 368 -78 374 78
rect 391 -78 397 78
rect 368 -103 397 -78
rect -397 -132 397 -103
<< mvpsubdiffcont >>
rect 374 -78 391 78
<< poly >>
rect -301 57 -251 65
rect -301 40 -293 57
rect -259 40 -251 57
rect -301 21 -251 40
rect -163 57 -113 65
rect -163 40 -155 57
rect -121 40 -113 57
rect -163 21 -113 40
rect -25 57 25 65
rect -25 40 -17 57
rect 17 40 25 57
rect -25 21 25 40
rect 113 57 163 65
rect 113 40 121 57
rect 155 40 163 57
rect 113 21 163 40
rect 251 57 301 65
rect 251 40 259 57
rect 293 40 301 57
rect 251 21 301 40
rect -301 -40 -251 -21
rect -301 -57 -293 -40
rect -259 -57 -251 -40
rect -301 -65 -251 -57
rect -163 -40 -113 -21
rect -163 -57 -155 -40
rect -121 -57 -113 -40
rect -163 -65 -113 -57
rect -25 -40 25 -21
rect -25 -57 -17 -40
rect 17 -57 25 -40
rect -25 -65 25 -57
rect 113 -40 163 -21
rect 113 -57 121 -40
rect 155 -57 163 -40
rect 113 -65 163 -57
rect 251 -40 301 -21
rect 251 -57 259 -40
rect 293 -57 301 -40
rect 251 -65 301 -57
<< polycont >>
rect -293 40 -259 57
rect -155 40 -121 57
rect -17 40 17 57
rect 121 40 155 57
rect 259 40 293 57
rect -293 -57 -259 -40
rect -155 -57 -121 -40
rect -17 -57 17 -40
rect 121 -57 155 -40
rect 259 -57 293 -40
<< locali >>
rect 374 78 391 86
rect -301 40 -293 57
rect -259 40 -251 57
rect -163 40 -155 57
rect -121 40 -113 57
rect -25 40 -17 57
rect 17 40 25 57
rect 113 40 121 57
rect 155 40 163 57
rect 251 40 259 57
rect 293 40 301 57
rect -324 15 -307 23
rect -324 -23 -307 -15
rect -245 15 -228 23
rect -245 -23 -228 -15
rect -186 15 -169 23
rect -186 -23 -169 -15
rect -107 15 -90 23
rect -107 -23 -90 -15
rect -48 15 -31 23
rect -48 -23 -31 -15
rect 31 15 48 23
rect 31 -23 48 -15
rect 90 15 107 23
rect 90 -23 107 -15
rect 169 15 186 23
rect 169 -23 186 -15
rect 228 15 245 23
rect 228 -23 245 -15
rect 307 15 324 23
rect 307 -23 324 -15
rect -301 -57 -293 -40
rect -259 -57 -251 -40
rect -163 -57 -155 -40
rect -121 -57 -113 -40
rect -25 -57 -17 -40
rect 17 -57 25 -40
rect 113 -57 121 -40
rect 155 -57 163 -40
rect 251 -57 259 -40
rect 293 -57 301 -40
rect 374 -86 391 -78
<< viali >>
rect -293 40 -259 57
rect -155 40 -121 57
rect -17 40 17 57
rect 121 40 155 57
rect 259 40 293 57
rect -324 -15 -307 15
rect -245 -15 -228 15
rect -186 -15 -169 15
rect -107 -15 -90 15
rect -48 -15 -31 15
rect 31 -15 48 15
rect 90 -15 107 15
rect 169 -15 186 15
rect 228 -15 245 15
rect 307 -15 324 15
rect -293 -57 -259 -40
rect -155 -57 -121 -40
rect -17 -57 17 -40
rect 121 -57 155 -40
rect 259 -57 293 -40
<< metal1 >>
rect -299 57 -253 60
rect -299 40 -293 57
rect -259 40 -253 57
rect -299 37 -253 40
rect -161 57 -115 60
rect -161 40 -155 57
rect -121 40 -115 57
rect -161 37 -115 40
rect -23 57 23 60
rect -23 40 -17 57
rect 17 40 23 57
rect -23 37 23 40
rect 115 57 161 60
rect 115 40 121 57
rect 155 40 161 57
rect 115 37 161 40
rect 253 57 299 60
rect 253 40 259 57
rect 293 40 299 57
rect 253 37 299 40
rect -327 15 -304 21
rect -327 -15 -324 15
rect -307 -15 -304 15
rect -327 -21 -304 -15
rect -248 15 -225 21
rect -248 -15 -245 15
rect -228 -15 -225 15
rect -248 -21 -225 -15
rect -189 15 -166 21
rect -189 -15 -186 15
rect -169 -15 -166 15
rect -189 -21 -166 -15
rect -110 15 -87 21
rect -110 -15 -107 15
rect -90 -15 -87 15
rect -110 -21 -87 -15
rect -51 15 -28 21
rect -51 -15 -48 15
rect -31 -15 -28 15
rect -51 -21 -28 -15
rect 28 15 51 21
rect 28 -15 31 15
rect 48 -15 51 15
rect 28 -21 51 -15
rect 87 15 110 21
rect 87 -15 90 15
rect 107 -15 110 15
rect 87 -21 110 -15
rect 166 15 189 21
rect 166 -15 169 15
rect 186 -15 189 15
rect 166 -21 189 -15
rect 225 15 248 21
rect 225 -15 228 15
rect 245 -15 248 15
rect 225 -21 248 -15
rect 304 15 327 21
rect 304 -15 307 15
rect 324 -15 327 15
rect 304 -21 327 -15
rect -299 -40 -253 -37
rect -299 -57 -293 -40
rect -259 -57 -253 -40
rect -299 -60 -253 -57
rect -161 -40 -115 -37
rect -161 -57 -155 -40
rect -121 -57 -115 -40
rect -161 -60 -115 -57
rect -23 -40 23 -37
rect -23 -57 -17 -40
rect 17 -57 23 -40
rect -23 -60 23 -57
rect 115 -40 161 -37
rect 115 -57 121 -40
rect 155 -57 161 -40
rect 115 -60 161 -57
rect 253 -40 299 -37
rect 253 -57 259 -40
rect 293 -57 299 -40
rect 253 -60 299 -57
<< properties >>
string FIXED_BBOX -382 -117 382 117
string gencell sky130_fd_pr__nfet_03v3_nvt
string library sky130
string parameters w 0.42 l 0.5 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 0 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
