magic
tech sky130A
magscale 1 2
timestamp 1717367797
<< pwell >>
rect 1152 -620 1232 -542
rect 1146 -846 1226 -768
<< locali >>
rect -274 -436 2605 -425
rect -274 -467 2606 -436
rect -274 -910 -232 -467
rect 46 -472 2606 -467
rect 46 -616 124 -472
rect 322 -618 400 -472
rect 600 -616 678 -472
rect 872 -616 950 -472
rect 1154 -616 1232 -574
rect 1426 -616 1504 -472
rect 1702 -618 1780 -472
rect 1976 -618 2054 -472
rect 2254 -616 2332 -472
rect 2528 -618 2606 -472
rect 50 -910 128 -774
rect 324 -910 402 -778
rect 600 -910 678 -778
rect 876 -910 954 -774
rect 1152 -816 1230 -774
rect 1424 -910 1502 -772
rect 1702 -910 1780 -774
rect 1980 -910 2058 -772
rect 2256 -910 2334 -772
rect 2532 -910 2610 -770
rect -274 -952 2612 -910
rect 690 -1090 806 -952
rect 690 -1134 712 -1090
rect 784 -1134 806 -1090
rect 690 -1160 806 -1134
rect 748 -1166 806 -1160
<< viali >>
rect 712 -1134 784 -1090
<< metal1 >>
rect 152 -428 3950 -374
rect -890 -790 -690 -590
rect -815 -990 -769 -790
rect -26 -990 6 -636
rect 158 -758 188 -428
rect 248 -758 278 -428
rect 440 -990 472 -634
rect 522 -990 554 -634
rect 710 -756 740 -428
rect 800 -758 830 -428
rect 1152 -552 1232 -542
rect 1152 -608 1154 -552
rect 1222 -608 1232 -552
rect 1152 -620 1232 -608
rect 992 -990 1024 -634
rect 1080 -990 1112 -636
rect 1264 -762 1294 -428
rect 1354 -764 1384 -428
rect 1146 -782 1226 -768
rect 1146 -838 1154 -782
rect 1222 -838 1226 -782
rect 1146 -846 1226 -838
rect 1540 -990 1572 -634
rect 1628 -990 1660 -636
rect 1814 -752 1844 -428
rect 1904 -752 1934 -428
rect 2092 -990 2124 -634
rect 2176 -990 2208 -642
rect 2368 -752 2398 -428
rect 2452 -750 2482 -428
rect 2642 -990 2674 -634
rect 2766 -848 2804 -428
rect 3893 -606 3947 -428
rect 3814 -806 4014 -606
rect -815 -1036 2678 -990
rect 2176 -1038 2208 -1036
rect 684 -1090 806 -1080
rect 684 -1134 712 -1090
rect 784 -1134 806 -1090
rect 684 -1316 806 -1134
rect 650 -1516 850 -1316
<< via1 >>
rect 1154 -608 1222 -552
rect 1154 -838 1222 -782
<< metal2 >>
rect 1146 -552 1232 -23
rect 1146 -608 1154 -552
rect 1222 -608 1232 -552
rect 1146 -616 1232 -608
rect 1146 -782 1232 -774
rect 1146 -838 1154 -782
rect 1222 -838 1232 -782
rect 1146 -1235 1232 -838
use sky130_fd_pr__nfet_03v3_nvt_J2JJF2  XM1
timestamp 1717366634
transform 1 0 1325 0 1 -695
box -1520 -300 1520 300
<< labels >>
flabel metal1 650 -1516 850 -1316 0 FreeSans 256 0 0 0 VG_H
port 0 nsew
flabel metal1 -890 -790 -690 -590 0 FreeSans 256 0 0 0 VD_H
port 1 nsew
flabel metal1 3814 -806 4014 -606 0 FreeSans 256 0 0 0 VLow_Src
port 2 nsew
<< end >>
