magic
tech sky130A
timestamp 1717363829
<< pwell >>
rect 500 -246 535 -187
rect 641 -245 676 -186
rect 499 -358 547 -322
rect 644 -358 675 -326
rect 757 -342 773 -260
rect 498 -379 675 -358
<< locali >>
rect -8 -192 676 -174
rect -8 -360 10 -192
rect 92 -245 127 -192
rect 226 -245 261 -192
rect 500 -246 535 -192
rect 641 -245 676 -192
rect 221 -360 268 -323
rect 499 -358 547 -322
rect 644 -358 675 -326
rect 498 -360 675 -358
rect -8 -361 675 -360
rect -8 -378 100 -361
rect 119 -378 675 -361
rect 498 -379 675 -378
<< viali >>
rect 100 -378 119 -361
<< metal1 >>
rect 336 352 425 438
rect 336 322 359 352
rect 406 322 425 352
rect 336 305 425 322
rect 357 201 408 205
rect 357 172 361 201
rect 404 172 408 201
rect 357 168 408 172
rect 0 -75 100 25
rect 675 -75 775 25
rect 49 -178 64 -75
rect 49 -192 624 -178
rect 49 -299 64 -192
rect 285 -313 302 -192
rect 324 -314 341 -192
rect 89 -361 123 -342
rect 89 -378 100 -361
rect 119 -378 123 -361
rect 89 -450 123 -378
rect 425 -396 444 -261
rect 462 -396 481 -262
rect 564 -313 581 -192
rect 599 -311 616 -192
rect 757 -261 774 -75
rect 697 -266 774 -261
rect 697 -296 773 -266
rect 757 -322 773 -296
rect 757 -396 775 -322
rect 425 -412 481 -396
rect 700 -412 775 -396
rect 75 -550 175 -450
rect 369 -607 420 -603
rect 369 -636 373 -607
rect 416 -636 420 -607
rect 369 -640 420 -636
rect 348 -771 437 -753
rect 348 -801 370 -771
rect 417 -801 437 -771
rect 348 -886 437 -801
<< via1 >>
rect 359 322 406 352
rect 361 172 404 201
rect 373 -636 416 -607
rect 370 -801 417 -771
<< metal2 >>
rect 339 352 425 362
rect 339 322 359 352
rect 406 322 425 352
rect 339 308 425 322
rect 357 201 408 308
rect 357 172 361 201
rect 404 172 408 201
rect 357 169 408 172
rect 369 -607 420 -605
rect 369 -636 373 -607
rect 416 -636 420 -607
rect 369 -759 420 -636
rect 349 -771 435 -759
rect 349 -801 370 -771
rect 417 -801 435 -771
rect 349 -813 435 -801
<< labels >>
flabel metal1 0 -75 100 25 0 FreeSans 128 0 0 0 VD_H
port 0 nsew
flabel metal1 75 -550 175 -450 0 FreeSans 128 0 0 0 VG_H
port 1 nsew
flabel metal1 675 -75 775 25 0 FreeSans 128 0 0 0 VLow_Src
port 2 nsew
<< end >>
