magic
tech sky130A
magscale 1 2
timestamp 1717277299
<< checkpaint >>
rect -1313 -2113 1629 4789
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
use sky130_fd_pr__nfet_01v8_ZJHFGD  XM3
timestamp 0
transform 1 0 158 0 1 1338
box -211 -2191 211 2191
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VD_H
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VG_H
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VLow_Src
port 2 nsew
<< end >>
