magic
tech sky130A
magscale 1 2
timestamp 1717370553
<< locali >>
rect 440 -928 538 -646
rect 712 -932 810 -650
rect 988 -936 1086 -654
rect 1266 -942 1364 -660
rect 1542 -946 1640 -664
rect 1816 -944 1914 -662
rect 2094 -946 2192 -664
rect 2372 -946 2470 -664
rect 2646 -946 2744 -664
rect 2924 -944 3022 -662
rect 3196 -936 3294 -654
rect 3472 -936 3570 -654
rect 3752 -942 3850 -660
rect 4020 -942 4118 -660
rect 4304 -946 4402 -664
rect 4578 -942 4676 -660
rect 4854 -946 4952 -664
rect 5128 -938 5226 -656
rect 5406 -946 5504 -664
rect 5676 -944 5774 -662
rect 5952 -938 6050 -656
rect 6234 -932 6332 -650
rect 6510 -936 6608 -654
rect 6784 -936 6882 -654
rect 7056 -936 7154 -654
rect 7338 -936 7436 -654
rect 7616 -942 7714 -660
rect 7890 -942 7988 -660
rect 8168 -946 8266 -664
rect 8444 -950 8542 -668
rect 8712 -950 8810 -668
rect 8994 -954 9092 -672
rect 9272 -952 9370 -670
rect 9546 -954 9644 -672
rect 9822 -954 9920 -672
rect 10092 -938 10190 -656
rect 10370 -946 10468 -664
rect 10652 -950 10750 -668
rect 10934 -946 11032 -664
rect 11202 -942 11300 -660
rect 11478 -942 11576 -660
rect 11748 -942 11846 -660
rect 12026 -936 12124 -654
rect 12308 -936 12406 -654
rect 12588 -936 12686 -654
rect 12854 -938 12952 -656
rect 13130 -944 13228 -662
rect 13410 -938 13508 -656
rect 13694 -938 13792 -656
rect 13972 -934 14070 -652
<< metal1 >>
rect -1366 -600 -1166 -400
rect 15478 -674 15678 -474
rect 4118 -1790 4318 -1590
use sky130_fd_pr__nfet_03v3_nvt_XW2EXC  XM1
timestamp 1717370147
transform 1 0 7113 0 1 -565
box -7178 -300 7178 300
<< labels >>
flabel metal1 4118 -1790 4318 -1590 0 FreeSans 256 0 0 0 VG_H
port 0 nsew
flabel metal1 -1366 -600 -1166 -400 0 FreeSans 256 0 0 0 VD_H
port 1 nsew
flabel metal1 15478 -674 15678 -474 0 FreeSans 256 0 0 0 VLow_Src
port 2 nsew
<< end >>
