magic
tech sky130A
magscale 1 2
timestamp 1717294976
<< error_p >>
rect -1310 -500 -1309 500
rect -1099 -500 -1098 500
rect -922 -500 -921 500
rect -711 -500 -710 500
rect 36 -500 37 500
rect 247 -500 248 500
rect 424 -500 425 500
rect 635 -500 636 500
rect 1382 -500 1383 500
rect 1593 -500 1594 500
<< nwell >>
rect -1784 -632 -1468 632
rect -552 -632 -122 632
rect 794 -632 1224 632
<< pwell >>
rect -2050 632 2050 898
rect -2050 -632 -1784 632
rect -1468 -632 -552 632
rect -122 -632 794 632
rect 1224 -632 2050 632
rect -2050 -898 2050 -632
<< mvnmos >>
rect -1309 -500 -1099 500
rect -921 -500 -711 500
rect 37 -500 247 500
rect 425 -500 635 500
rect 1383 -500 1593 500
<< mvndiff >>
rect -1099 488 -1041 500
rect -1099 -488 -1087 488
rect -1053 -488 -1041 488
rect -1099 -500 -1041 -488
rect -979 488 -921 500
rect -979 -488 -967 488
rect -933 -488 -921 488
rect -979 -500 -921 -488
rect 247 488 305 500
rect 247 -488 259 488
rect 293 -488 305 488
rect 247 -500 305 -488
rect 367 488 425 500
rect 367 -488 379 488
rect 413 -488 425 488
rect 367 -500 425 -488
rect 1593 488 1651 500
rect 1593 -488 1605 488
rect 1639 -488 1651 488
rect 1593 -500 1651 -488
<< mvndiffc >>
rect -1087 -488 -1053 488
rect -967 -488 -933 488
rect 259 -488 293 488
rect 379 -488 413 488
rect 1605 -488 1639 488
<< mvpsubdiff >>
rect -2014 850 2014 862
rect -2014 816 -1906 850
rect 1906 816 2014 850
rect -2014 804 2014 816
rect -2014 754 -1956 804
rect -2014 -754 -2002 754
rect -1968 -754 -1956 754
rect 1956 754 2014 804
rect -2014 -804 -1956 -754
rect 1956 -754 1968 754
rect 2002 -754 2014 754
rect 1956 -804 2014 -754
rect -2014 -816 2014 -804
rect -2014 -850 -1906 -816
rect 1906 -850 2014 -816
rect -2014 -862 2014 -850
<< mvnsubdiff >>
rect -1652 476 -1600 500
rect -1652 -476 -1643 476
rect -1609 -476 -1600 476
rect -1652 -500 -1600 -476
rect -420 476 -368 500
rect -420 -476 -411 476
rect -377 -476 -368 476
rect -420 -500 -368 -476
rect -306 476 -254 500
rect -306 -476 -297 476
rect -263 -476 -254 476
rect -306 -500 -254 -476
rect 926 476 978 500
rect 926 -476 935 476
rect 969 -476 978 476
rect 926 -500 978 -476
rect 1040 476 1092 500
rect 1040 -476 1049 476
rect 1083 -476 1092 476
rect 1040 -500 1092 -476
<< mvpsubdiffcont >>
rect -1906 816 1906 850
rect -2002 -754 -1968 754
rect 1968 -754 2002 754
rect -1906 -850 1906 -816
<< mvnsubdiffcont >>
rect -1643 -476 -1609 476
rect -411 -476 -377 476
rect -297 -476 -263 476
rect 935 -476 969 476
rect 1049 -476 1083 476
<< extdrain >>
rect -1600 -500 -1309 500
rect -711 -500 -420 500
rect -254 -500 37 500
rect 635 -500 926 500
rect 1092 -500 1383 500
<< poly >>
rect -1309 572 -1099 588
rect -1309 538 -1293 572
rect -1115 538 -1099 572
rect -1309 500 -1099 538
rect -921 572 -711 588
rect -921 538 -905 572
rect -727 538 -711 572
rect -921 500 -711 538
rect 37 572 247 588
rect 37 538 53 572
rect 231 538 247 572
rect 37 500 247 538
rect 425 572 635 588
rect 425 538 441 572
rect 619 538 635 572
rect 425 500 635 538
rect 1383 572 1593 588
rect 1383 538 1399 572
rect 1577 538 1593 572
rect 1383 500 1593 538
rect -1309 -538 -1099 -500
rect -1309 -572 -1293 -538
rect -1115 -572 -1099 -538
rect -1309 -588 -1099 -572
rect -921 -538 -711 -500
rect -921 -572 -905 -538
rect -727 -572 -711 -538
rect -921 -588 -711 -572
rect 37 -538 247 -500
rect 37 -572 53 -538
rect 231 -572 247 -538
rect 37 -588 247 -572
rect 425 -538 635 -500
rect 425 -572 441 -538
rect 619 -572 635 -538
rect 425 -588 635 -572
rect 1383 -538 1593 -500
rect 1383 -572 1399 -538
rect 1577 -572 1593 -538
rect 1383 -588 1593 -572
<< polycont >>
rect -1293 538 -1115 572
rect -905 538 -727 572
rect 53 538 231 572
rect 441 538 619 572
rect 1399 538 1577 572
rect -1293 -572 -1115 -538
rect -905 -572 -727 -538
rect 53 -572 231 -538
rect 441 -572 619 -538
rect 1399 -572 1577 -538
<< locali >>
rect -2002 816 -1906 850
rect 1906 816 2002 850
rect -2002 754 -1968 816
rect 1968 754 2002 816
rect -1309 538 -1293 572
rect -1115 538 -1099 572
rect -921 538 -905 572
rect -727 538 -711 572
rect 37 538 53 572
rect 231 538 247 572
rect 425 538 441 572
rect 619 538 635 572
rect 1383 538 1399 572
rect 1577 538 1593 572
rect -1643 488 -1609 492
rect -1643 -492 -1609 -488
rect -1087 488 -1053 504
rect -1087 -504 -1053 -488
rect -967 488 -933 504
rect -967 -504 -933 -488
rect -411 488 -377 492
rect -411 -492 -377 -488
rect -297 488 -263 492
rect -297 -492 -263 -488
rect 259 488 293 504
rect 259 -504 293 -488
rect 379 488 413 504
rect 379 -504 413 -488
rect 935 488 969 492
rect 935 -492 969 -488
rect 1049 488 1083 492
rect 1049 -492 1083 -488
rect 1605 488 1639 504
rect 1605 -504 1639 -488
rect -1309 -572 -1293 -538
rect -1115 -572 -1099 -538
rect -921 -572 -905 -538
rect -727 -572 -711 -538
rect 37 -572 53 -538
rect 231 -572 247 -538
rect 425 -572 441 -538
rect 619 -572 635 -538
rect 1383 -572 1399 -538
rect 1577 -572 1593 -538
rect -2002 -816 -1968 -754
rect 1968 -816 2002 -754
rect -2002 -850 -1906 -816
rect 1906 -850 2002 -816
<< viali >>
rect -1293 538 -1115 572
rect -905 538 -727 572
rect 53 538 231 572
rect 441 538 619 572
rect 1399 538 1577 572
rect -1643 476 -1609 488
rect -1643 -476 -1609 476
rect -1643 -488 -1609 -476
rect -1087 -488 -1053 488
rect -967 -488 -933 488
rect -411 476 -377 488
rect -411 -476 -377 476
rect -411 -488 -377 -476
rect -297 476 -263 488
rect -297 -476 -263 476
rect -297 -488 -263 -476
rect 259 -488 293 488
rect 379 -488 413 488
rect 935 476 969 488
rect 935 -476 969 476
rect 935 -488 969 -476
rect 1049 476 1083 488
rect 1049 -476 1083 476
rect 1049 -488 1083 -476
rect 1605 -488 1639 488
rect -1293 -572 -1115 -538
rect -905 -572 -727 -538
rect 53 -572 231 -538
rect 441 -572 619 -538
rect 1399 -572 1577 -538
<< metal1 >>
rect -1305 572 -1103 578
rect -1305 538 -1293 572
rect -1115 538 -1103 572
rect -1305 532 -1103 538
rect -917 572 -715 578
rect -917 538 -905 572
rect -727 538 -715 572
rect -917 532 -715 538
rect 41 572 243 578
rect 41 538 53 572
rect 231 538 243 572
rect 41 532 243 538
rect 429 572 631 578
rect 429 538 441 572
rect 619 538 631 572
rect 429 532 631 538
rect 1387 572 1589 578
rect 1387 538 1399 572
rect 1577 538 1589 572
rect 1387 532 1589 538
rect -1649 488 -1603 500
rect -1649 -488 -1643 488
rect -1609 -488 -1603 488
rect -1649 -500 -1603 -488
rect -1093 488 -1047 500
rect -1093 -488 -1087 488
rect -1053 -488 -1047 488
rect -1093 -500 -1047 -488
rect -973 488 -927 500
rect -973 -488 -967 488
rect -933 -488 -927 488
rect -973 -500 -927 -488
rect -417 488 -371 500
rect -417 -488 -411 488
rect -377 -488 -371 488
rect -417 -500 -371 -488
rect -303 488 -257 500
rect -303 -488 -297 488
rect -263 -488 -257 488
rect -303 -500 -257 -488
rect 253 488 299 500
rect 253 -488 259 488
rect 293 -488 299 488
rect 253 -500 299 -488
rect 373 488 419 500
rect 373 -488 379 488
rect 413 -488 419 488
rect 373 -500 419 -488
rect 929 488 975 500
rect 929 -488 935 488
rect 969 -488 975 488
rect 929 -500 975 -488
rect 1043 488 1089 500
rect 1043 -488 1049 488
rect 1083 -488 1089 488
rect 1043 -500 1089 -488
rect 1599 488 1645 500
rect 1599 -488 1605 488
rect 1639 -488 1645 488
rect 1599 -500 1645 -488
rect -1305 -538 -1103 -532
rect -1305 -572 -1293 -538
rect -1115 -572 -1103 -538
rect -1305 -578 -1103 -572
rect -917 -538 -715 -532
rect -917 -572 -905 -538
rect -727 -572 -715 -538
rect -917 -578 -715 -572
rect 41 -538 243 -532
rect 41 -572 53 -538
rect 231 -572 243 -538
rect 41 -578 243 -572
rect 429 -538 631 -532
rect 429 -572 441 -538
rect 619 -572 631 -538
rect 429 -578 631 -572
rect 1387 -538 1589 -532
rect 1387 -572 1399 -538
rect 1577 -572 1589 -538
rect 1387 -578 1589 -572
<< properties >>
string FIXED_BBOX -1985 -833 1985 833
string gencell sky130_fd_pr__nfet_g5v0d16v0
string library sky130
string parameters w 5.00 l 1.050 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 1.050 wmin 5.00 full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
