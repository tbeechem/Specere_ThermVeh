magic
tech sky130A
timestamp 1717702195
use GSense_Contacts_nFET_3V_1nf  GSense_Contacts_nFET_3V_1nf_0
timestamp 1717698305
transform 1 0 209100 0 1 28982
box -14400 -14282 15900 13218
use GSense_Contacts_nFET_3V_1nf  GSense_Contacts_nFET_3V_1nf_1
timestamp 1717698305
transform 1 0 74100 0 1 28982
box -14400 -14282 15900 13218
use GSense_Contacts_nFET_3V_1nf  GSense_Contacts_nFET_3V_1nf_2
timestamp 1717698305
transform 1 0 29100 0 1 291482
box -14400 -14282 15900 13218
use GSense_Contacts_nFET_3V_1nf  GSense_Contacts_nFET_3V_1nf_3
timestamp 1717698305
transform 1 0 29100 0 1 328982
box -14400 -14282 15900 13218
use GSense_Contacts_nFT_g5_10Vd_1nf  GSense_Contacts_nFT_g5_10Vd_1nf_0
timestamp 1717698512
transform 1 0 119100 0 1 28982
box -14400 -14282 15800 13318
use GSense_Contacts_nFT_g5_10Vd_1nf  GSense_Contacts_nFT_g5_10Vd_1nf_1
timestamp 1717698512
transform 1 0 254100 0 1 28982
box -14400 -14282 15800 13318
use GSense_Contacts_nFT_g5_10Vd_1nf  GSense_Contacts_nFT_g5_10Vd_1nf_2
timestamp 1717698512
transform 1 0 74100 0 1 291482
box -14400 -14282 15800 13318
use GSense_Contacts_pfet_1p8Vd_1p8Vg  GSense_Contacts_pfet_1p8Vd_1p8Vg_0
timestamp 1717699159
transform 1 0 29100 0 1 73982
box -14399 -14220 16001 13180
use GSense_Contacts_pfet_1p8Vd_1p8Vg  GSense_Contacts_pfet_1p8Vd_1p8Vg_1
timestamp 1717699159
transform 1 0 164100 0 1 73982
box -14399 -14220 16001 13180
use GSense_Contacts_pfet_1p8Vd_1p8Vg  GSense_Contacts_pfet_1p8Vd_1p8Vg_2
timestamp 1717699159
transform 1 0 119100 0 1 328982
box -14399 -14220 16001 13180
use GSense_nFET_1W015L_1F_Contacts  GSense_nFET_1W015L_1F_Contacts_0
timestamp 1717698710
transform 1 0 119100 0 1 73982
box -14300 -14282 15900 13218
use GSense_nFET_1W015L_1F_Contacts  GSense_nFET_1W015L_1F_Contacts_1
timestamp 1717698710
transform 1 0 164100 0 1 28982
box -14300 -14282 15900 13218
use GSense_nFET_1W015L_1F_Contacts  GSense_nFET_1W015L_1F_Contacts_2
timestamp 1717698710
transform 1 0 29100 0 1 28982
box -14300 -14282 15900 13218
use GSense_nFET_1W015L_1F_Contacts  GSense_nFET_1W015L_1F_Contacts_3
timestamp 1717698710
transform 1 0 254100 0 1 73982
box -14300 -14282 15900 13218
use GSense_nFET_1W015L_1F_Contacts  GSense_nFET_1W015L_1F_Contacts_4
timestamp 1717698710
transform 1 0 119100 0 1 291482
box -14300 -14282 15900 13218
use GSense_nFET_1W015L_1F_Contacts  GSense_nFET_1W015L_1F_Contacts_5
timestamp 1717698710
transform 1 0 74100 0 1 328982
box -14300 -14282 15900 13218
use GSense_nFET_3p3V_5nF_Contacts_V2  GSense_nFET_3p3V_5nF_Contacts_V2_0
timestamp 1717699633
transform 1 0 29100 0 1 127032
box -14299 -22370 15901 21330
use GSense_nFET_3p3V_5nF_Contacts_V2  GSense_nFET_3p3V_5nF_Contacts_V2_1
timestamp 1717699633
transform 1 0 254100 0 1 187032
box -14299 -22370 15901 21330
use GSense_nFET_3p3V_5nF_Contacts_V2  GSense_nFET_3p3V_5nF_Contacts_V2_2
timestamp 1717699633
transform 1 0 209100 0 1 247032
box -14299 -22370 15901 21330
use GSense_pFET_10Vd_5p5Vg_1nf  GSense_pFET_10Vd_5p5Vg_1nf_0
timestamp 1717698855
transform 1 0 74100 0 1 73982
box -14400 -14282 15800 13218
use GSense_pFET_10Vd_5p5Vg_1nf  GSense_pFET_10Vd_5p5Vg_1nf_1
timestamp 1717698855
transform 1 0 209100 0 1 73982
box -14400 -14282 15800 13218
use GSense_pFET_10Vd_5p5Vg_1nf  GSense_pFET_10Vd_5p5Vg_1nf_2
timestamp 1717698855
transform 1 0 164100 0 1 291482
box -14400 -14282 15800 13218
use nFET_3p3Vd_3VG_51NF_LTherm_Contacts  nFET_3p3Vd_3VG_51NF_LTherm_Contacts_0
timestamp 1717699946
transform 1 0 119289 0 1 126836
box -14388 -22374 15912 21426
use nFET_3p3Vd_3VG_51NF_LTherm_Contacts  nFET_3p3Vd_3VG_51NF_LTherm_Contacts_1
timestamp 1717699946
transform 1 0 164100 0 1 247032
box -14388 -22374 15912 21426
use nFET_3p3Vd_3VG_51NF_LTherm_Contacts  nFET_3p3Vd_3VG_51NF_LTherm_Contacts_2
timestamp 1717699946
transform 1 0 164100 0 1 187032
box -14388 -22374 15912 21426
use nFET_3VD_3VG_10nF_Contacts  nFET_3VD_3VG_10nF_Contacts_0
timestamp 1717699946
transform 1 0 73662 0 1 126930
box -14361 -22368 15839 21432
use nFET_3VD_3VG_10nF_Contacts  nFET_3VD_3VG_10nF_Contacts_1
timestamp 1717699946
transform 1 0 254100 0 1 247032
box -14361 -22368 15839 21432
use nFET_3VD_3VG_10nF_Contacts  nFET_3VD_3VG_10nF_Contacts_2
timestamp 1717699946
transform 1 0 209100 0 1 187032
box -14361 -22368 15839 21432
use nFET_3VD_3VG_10nF_Contacts  nFET_3VD_3VG_10nF_Contacts_3
timestamp 1717699946
transform 1 0 29100 0 1 247032
box -14361 -22368 15839 21432
use nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts  nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_0
timestamp 1717702195
transform 1 0 209100 0 1 127032
box -14399 -22370 15901 21430
use nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts  nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_1
timestamp 1717702195
transform 1 0 254100 0 1 127032
box -14399 -22370 15901 21430
use nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts  nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_2
timestamp 1717702195
transform 1 0 29100 0 1 187032
box -14399 -22370 15901 21430
use nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts  nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_3
timestamp 1717702195
transform 1 0 74100 0 1 247032
box -14399 -22370 15901 21430
use nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts  nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_5
timestamp 1717702195
transform 1 0 74100 0 1 187032
box -14399 -22370 15901 21430
use nFET_3VD_3VG_50nF_Therm_FET12  nFET_3VD_3VG_50nF_Therm_FET12_0
timestamp 1717700119
transform 1 0 164100 0 1 127032
box -14399 -22370 15901 21230
use nFET_3VD_3VG_50nF_Therm_FET12  nFET_3VD_3VG_50nF_Therm_FET12_1
timestamp 1717700119
transform 1 0 119100 0 1 247032
box -14399 -22370 15901 21230
use nFET_3VD_3VG_50nF_Therm_FET12  nFET_3VD_3VG_50nF_Therm_FET12_3
timestamp 1717700119
transform 1 0 119100 0 1 187032
box -14399 -22370 15901 21230
<< end >>
