magic
tech sky130A
magscale 1 2
timestamp 1717469809
<< nwell >>
rect 419065 656969 419681 657763
rect 239145 655527 239567 656165
rect 329263 580045 329879 580839
rect 59145 145527 59567 146165
rect 149263 145045 149879 145839
rect 329145 145527 329567 146165
rect 419263 145045 419879 145839
<< pwell >>
rect 328964 657498 329386 658118
rect 508964 657498 509386 658118
rect 59383 655525 59939 656241
rect 149162 655574 149584 656194
rect 419185 582449 419741 583165
rect 509195 582159 509751 582875
rect 59383 580525 59939 581241
rect 149393 580235 149949 580951
rect 239162 580574 239584 581194
rect 337132 492417 337230 492480
rect 337402 492417 337500 492478
rect 58659 491429 61699 492029
rect 323649 491817 338005 492417
rect 156592 491739 156690 491803
rect 156862 491739 156960 491801
rect 143109 491139 157465 491739
rect 245949 491143 246047 491207
rect 246219 491143 246317 491205
rect 232466 490543 246822 491143
rect 418658 491101 420318 491701
rect 508659 491429 511699 492029
rect 337132 372417 337230 372480
rect 337402 372417 337500 372478
rect 323649 371817 338005 372417
rect 66592 371739 66690 371803
rect 66862 371739 66960 371801
rect 156592 371739 156690 371803
rect 156862 371739 156960 371801
rect 53109 371139 67465 371739
rect 143109 371139 157465 371739
rect 418659 371429 421699 372029
rect 245949 371143 246047 371207
rect 246219 371143 246317 371205
rect 232466 370543 246822 371143
rect 508658 371101 510318 371701
rect 247510 252025 247608 252088
rect 247780 252025 247878 252086
rect 58658 251101 60318 251701
rect 147783 251225 150823 251825
rect 234027 251425 248383 252025
rect 426592 251739 426690 251803
rect 426862 251739 426960 251801
rect 516592 251739 516690 251803
rect 516862 251739 516960 251801
rect 335949 251143 336047 251207
rect 336219 251143 336317 251205
rect 322466 250543 336822 251143
rect 413109 251139 427465 251739
rect 503109 251139 517465 251739
rect 239162 145574 239584 146194
rect 509162 145574 509584 146194
rect 59162 55574 59584 56194
rect 149383 55525 149939 56241
rect 239393 55235 239949 55951
rect 329162 55574 329584 56194
rect 419383 55525 419939 56241
rect 509393 55235 509949 55951
<< nmos >>
rect 329160 657708 329190 657908
rect 509160 657708 509190 657908
rect 149358 655784 149388 655984
rect 239358 580784 239388 580984
rect 239358 145784 239388 145984
rect 509358 145784 509388 145984
rect 59358 55784 59388 55984
rect 329358 55784 329388 55984
<< pmos >>
rect 239341 655746 239371 655946
rect 59341 145746 59371 145946
rect 329341 145746 329371 145946
<< nnmos >>
rect 59611 655783 59711 655983
rect 419413 582707 419513 582907
rect 59611 580783 59711 580983
rect 58887 491687 58987 491771
rect 59163 491687 59263 491771
rect 59439 491687 59539 491771
rect 59715 491687 59815 491771
rect 59991 491687 60091 491771
rect 60267 491687 60367 491771
rect 60543 491687 60643 491771
rect 60819 491687 60919 491771
rect 61095 491687 61195 491771
rect 61371 491687 61471 491771
rect 323877 492075 323977 492159
rect 324153 492075 324253 492159
rect 324429 492075 324529 492159
rect 324705 492075 324805 492159
rect 324981 492075 325081 492159
rect 325257 492075 325357 492159
rect 325533 492075 325633 492159
rect 325809 492075 325909 492159
rect 326085 492075 326185 492159
rect 326361 492075 326461 492159
rect 326637 492075 326737 492159
rect 326913 492075 327013 492159
rect 327189 492075 327289 492159
rect 327465 492075 327565 492159
rect 327741 492075 327841 492159
rect 328017 492075 328117 492159
rect 328293 492075 328393 492159
rect 328569 492075 328669 492159
rect 328845 492075 328945 492159
rect 329121 492075 329221 492159
rect 329397 492075 329497 492159
rect 329673 492075 329773 492159
rect 329949 492075 330049 492159
rect 330225 492075 330325 492159
rect 330501 492075 330601 492159
rect 330777 492075 330877 492159
rect 331053 492075 331153 492159
rect 331329 492075 331429 492159
rect 331605 492075 331705 492159
rect 331881 492075 331981 492159
rect 332157 492075 332257 492159
rect 332433 492075 332533 492159
rect 332709 492075 332809 492159
rect 332985 492075 333085 492159
rect 333261 492075 333361 492159
rect 333537 492075 333637 492159
rect 333813 492075 333913 492159
rect 334089 492075 334189 492159
rect 334365 492075 334465 492159
rect 334641 492075 334741 492159
rect 334917 492075 335017 492159
rect 335193 492075 335293 492159
rect 335469 492075 335569 492159
rect 335745 492075 335845 492159
rect 336021 492075 336121 492159
rect 336297 492075 336397 492159
rect 336573 492075 336673 492159
rect 336849 492075 336949 492159
rect 337125 492075 337225 492159
rect 337401 492075 337501 492159
rect 337677 492075 337777 492159
rect 143337 491397 143437 491481
rect 143613 491397 143713 491481
rect 143889 491397 143989 491481
rect 144165 491397 144265 491481
rect 144441 491397 144541 491481
rect 144717 491397 144817 491481
rect 144993 491397 145093 491481
rect 145269 491397 145369 491481
rect 145545 491397 145645 491481
rect 145821 491397 145921 491481
rect 146097 491397 146197 491481
rect 146373 491397 146473 491481
rect 146649 491397 146749 491481
rect 146925 491397 147025 491481
rect 147201 491397 147301 491481
rect 147477 491397 147577 491481
rect 147753 491397 147853 491481
rect 148029 491397 148129 491481
rect 148305 491397 148405 491481
rect 148581 491397 148681 491481
rect 148857 491397 148957 491481
rect 149133 491397 149233 491481
rect 149409 491397 149509 491481
rect 149685 491397 149785 491481
rect 149961 491397 150061 491481
rect 150237 491397 150337 491481
rect 150513 491397 150613 491481
rect 150789 491397 150889 491481
rect 151065 491397 151165 491481
rect 151341 491397 151441 491481
rect 151617 491397 151717 491481
rect 151893 491397 151993 491481
rect 152169 491397 152269 491481
rect 152445 491397 152545 491481
rect 152721 491397 152821 491481
rect 152997 491397 153097 491481
rect 153273 491397 153373 491481
rect 153549 491397 153649 491481
rect 153825 491397 153925 491481
rect 154101 491397 154201 491481
rect 154377 491397 154477 491481
rect 154653 491397 154753 491481
rect 154929 491397 155029 491481
rect 155205 491397 155305 491481
rect 155481 491397 155581 491481
rect 155757 491397 155857 491481
rect 156033 491397 156133 491481
rect 156309 491397 156409 491481
rect 156585 491397 156685 491481
rect 156861 491397 156961 491481
rect 157137 491397 157237 491481
rect 418886 491359 418986 491443
rect 419162 491359 419262 491443
rect 419438 491359 419538 491443
rect 419714 491359 419814 491443
rect 419990 491359 420090 491443
rect 508887 491687 508987 491771
rect 509163 491687 509263 491771
rect 509439 491687 509539 491771
rect 509715 491687 509815 491771
rect 509991 491687 510091 491771
rect 510267 491687 510367 491771
rect 510543 491687 510643 491771
rect 510819 491687 510919 491771
rect 511095 491687 511195 491771
rect 511371 491687 511471 491771
rect 232694 490801 232794 490885
rect 232970 490801 233070 490885
rect 233246 490801 233346 490885
rect 233522 490801 233622 490885
rect 233798 490801 233898 490885
rect 234074 490801 234174 490885
rect 234350 490801 234450 490885
rect 234626 490801 234726 490885
rect 234902 490801 235002 490885
rect 235178 490801 235278 490885
rect 235454 490801 235554 490885
rect 235730 490801 235830 490885
rect 236006 490801 236106 490885
rect 236282 490801 236382 490885
rect 236558 490801 236658 490885
rect 236834 490801 236934 490885
rect 237110 490801 237210 490885
rect 237386 490801 237486 490885
rect 237662 490801 237762 490885
rect 237938 490801 238038 490885
rect 238214 490801 238314 490885
rect 238490 490801 238590 490885
rect 238766 490801 238866 490885
rect 239042 490801 239142 490885
rect 239318 490801 239418 490885
rect 239594 490801 239694 490885
rect 239870 490801 239970 490885
rect 240146 490801 240246 490885
rect 240422 490801 240522 490885
rect 240698 490801 240798 490885
rect 240974 490801 241074 490885
rect 241250 490801 241350 490885
rect 241526 490801 241626 490885
rect 241802 490801 241902 490885
rect 242078 490801 242178 490885
rect 242354 490801 242454 490885
rect 242630 490801 242730 490885
rect 242906 490801 243006 490885
rect 243182 490801 243282 490885
rect 243458 490801 243558 490885
rect 243734 490801 243834 490885
rect 244010 490801 244110 490885
rect 244286 490801 244386 490885
rect 244562 490801 244662 490885
rect 244838 490801 244938 490885
rect 245114 490801 245214 490885
rect 245390 490801 245490 490885
rect 245666 490801 245766 490885
rect 245942 490801 246042 490885
rect 246218 490801 246318 490885
rect 246494 490801 246594 490885
rect 323877 372075 323977 372159
rect 324153 372075 324253 372159
rect 324429 372075 324529 372159
rect 324705 372075 324805 372159
rect 324981 372075 325081 372159
rect 325257 372075 325357 372159
rect 325533 372075 325633 372159
rect 325809 372075 325909 372159
rect 326085 372075 326185 372159
rect 326361 372075 326461 372159
rect 326637 372075 326737 372159
rect 326913 372075 327013 372159
rect 327189 372075 327289 372159
rect 327465 372075 327565 372159
rect 327741 372075 327841 372159
rect 328017 372075 328117 372159
rect 328293 372075 328393 372159
rect 328569 372075 328669 372159
rect 328845 372075 328945 372159
rect 329121 372075 329221 372159
rect 329397 372075 329497 372159
rect 329673 372075 329773 372159
rect 329949 372075 330049 372159
rect 330225 372075 330325 372159
rect 330501 372075 330601 372159
rect 330777 372075 330877 372159
rect 331053 372075 331153 372159
rect 331329 372075 331429 372159
rect 331605 372075 331705 372159
rect 331881 372075 331981 372159
rect 332157 372075 332257 372159
rect 332433 372075 332533 372159
rect 332709 372075 332809 372159
rect 332985 372075 333085 372159
rect 333261 372075 333361 372159
rect 333537 372075 333637 372159
rect 333813 372075 333913 372159
rect 334089 372075 334189 372159
rect 334365 372075 334465 372159
rect 334641 372075 334741 372159
rect 334917 372075 335017 372159
rect 335193 372075 335293 372159
rect 335469 372075 335569 372159
rect 335745 372075 335845 372159
rect 336021 372075 336121 372159
rect 336297 372075 336397 372159
rect 336573 372075 336673 372159
rect 336849 372075 336949 372159
rect 337125 372075 337225 372159
rect 337401 372075 337501 372159
rect 337677 372075 337777 372159
rect 53337 371397 53437 371481
rect 53613 371397 53713 371481
rect 53889 371397 53989 371481
rect 54165 371397 54265 371481
rect 54441 371397 54541 371481
rect 54717 371397 54817 371481
rect 54993 371397 55093 371481
rect 55269 371397 55369 371481
rect 55545 371397 55645 371481
rect 55821 371397 55921 371481
rect 56097 371397 56197 371481
rect 56373 371397 56473 371481
rect 56649 371397 56749 371481
rect 56925 371397 57025 371481
rect 57201 371397 57301 371481
rect 57477 371397 57577 371481
rect 57753 371397 57853 371481
rect 58029 371397 58129 371481
rect 58305 371397 58405 371481
rect 58581 371397 58681 371481
rect 58857 371397 58957 371481
rect 59133 371397 59233 371481
rect 59409 371397 59509 371481
rect 59685 371397 59785 371481
rect 59961 371397 60061 371481
rect 60237 371397 60337 371481
rect 60513 371397 60613 371481
rect 60789 371397 60889 371481
rect 61065 371397 61165 371481
rect 61341 371397 61441 371481
rect 61617 371397 61717 371481
rect 61893 371397 61993 371481
rect 62169 371397 62269 371481
rect 62445 371397 62545 371481
rect 62721 371397 62821 371481
rect 62997 371397 63097 371481
rect 63273 371397 63373 371481
rect 63549 371397 63649 371481
rect 63825 371397 63925 371481
rect 64101 371397 64201 371481
rect 64377 371397 64477 371481
rect 64653 371397 64753 371481
rect 64929 371397 65029 371481
rect 65205 371397 65305 371481
rect 65481 371397 65581 371481
rect 65757 371397 65857 371481
rect 66033 371397 66133 371481
rect 66309 371397 66409 371481
rect 66585 371397 66685 371481
rect 66861 371397 66961 371481
rect 67137 371397 67237 371481
rect 143337 371397 143437 371481
rect 143613 371397 143713 371481
rect 143889 371397 143989 371481
rect 144165 371397 144265 371481
rect 144441 371397 144541 371481
rect 144717 371397 144817 371481
rect 144993 371397 145093 371481
rect 145269 371397 145369 371481
rect 145545 371397 145645 371481
rect 145821 371397 145921 371481
rect 146097 371397 146197 371481
rect 146373 371397 146473 371481
rect 146649 371397 146749 371481
rect 146925 371397 147025 371481
rect 147201 371397 147301 371481
rect 147477 371397 147577 371481
rect 147753 371397 147853 371481
rect 148029 371397 148129 371481
rect 148305 371397 148405 371481
rect 148581 371397 148681 371481
rect 148857 371397 148957 371481
rect 149133 371397 149233 371481
rect 149409 371397 149509 371481
rect 149685 371397 149785 371481
rect 149961 371397 150061 371481
rect 150237 371397 150337 371481
rect 150513 371397 150613 371481
rect 150789 371397 150889 371481
rect 151065 371397 151165 371481
rect 151341 371397 151441 371481
rect 151617 371397 151717 371481
rect 151893 371397 151993 371481
rect 152169 371397 152269 371481
rect 152445 371397 152545 371481
rect 152721 371397 152821 371481
rect 152997 371397 153097 371481
rect 153273 371397 153373 371481
rect 153549 371397 153649 371481
rect 153825 371397 153925 371481
rect 154101 371397 154201 371481
rect 154377 371397 154477 371481
rect 154653 371397 154753 371481
rect 154929 371397 155029 371481
rect 155205 371397 155305 371481
rect 155481 371397 155581 371481
rect 155757 371397 155857 371481
rect 156033 371397 156133 371481
rect 156309 371397 156409 371481
rect 156585 371397 156685 371481
rect 156861 371397 156961 371481
rect 157137 371397 157237 371481
rect 418887 371687 418987 371771
rect 419163 371687 419263 371771
rect 419439 371687 419539 371771
rect 419715 371687 419815 371771
rect 419991 371687 420091 371771
rect 420267 371687 420367 371771
rect 420543 371687 420643 371771
rect 420819 371687 420919 371771
rect 421095 371687 421195 371771
rect 421371 371687 421471 371771
rect 508886 371359 508986 371443
rect 509162 371359 509262 371443
rect 509438 371359 509538 371443
rect 509714 371359 509814 371443
rect 509990 371359 510090 371443
rect 232694 370801 232794 370885
rect 232970 370801 233070 370885
rect 233246 370801 233346 370885
rect 233522 370801 233622 370885
rect 233798 370801 233898 370885
rect 234074 370801 234174 370885
rect 234350 370801 234450 370885
rect 234626 370801 234726 370885
rect 234902 370801 235002 370885
rect 235178 370801 235278 370885
rect 235454 370801 235554 370885
rect 235730 370801 235830 370885
rect 236006 370801 236106 370885
rect 236282 370801 236382 370885
rect 236558 370801 236658 370885
rect 236834 370801 236934 370885
rect 237110 370801 237210 370885
rect 237386 370801 237486 370885
rect 237662 370801 237762 370885
rect 237938 370801 238038 370885
rect 238214 370801 238314 370885
rect 238490 370801 238590 370885
rect 238766 370801 238866 370885
rect 239042 370801 239142 370885
rect 239318 370801 239418 370885
rect 239594 370801 239694 370885
rect 239870 370801 239970 370885
rect 240146 370801 240246 370885
rect 240422 370801 240522 370885
rect 240698 370801 240798 370885
rect 240974 370801 241074 370885
rect 241250 370801 241350 370885
rect 241526 370801 241626 370885
rect 241802 370801 241902 370885
rect 242078 370801 242178 370885
rect 242354 370801 242454 370885
rect 242630 370801 242730 370885
rect 242906 370801 243006 370885
rect 243182 370801 243282 370885
rect 243458 370801 243558 370885
rect 243734 370801 243834 370885
rect 244010 370801 244110 370885
rect 244286 370801 244386 370885
rect 244562 370801 244662 370885
rect 244838 370801 244938 370885
rect 245114 370801 245214 370885
rect 245390 370801 245490 370885
rect 245666 370801 245766 370885
rect 245942 370801 246042 370885
rect 246218 370801 246318 370885
rect 246494 370801 246594 370885
rect 58886 251359 58986 251443
rect 59162 251359 59262 251443
rect 59438 251359 59538 251443
rect 59714 251359 59814 251443
rect 59990 251359 60090 251443
rect 148011 251483 148111 251567
rect 148287 251483 148387 251567
rect 148563 251483 148663 251567
rect 148839 251483 148939 251567
rect 149115 251483 149215 251567
rect 149391 251483 149491 251567
rect 149667 251483 149767 251567
rect 149943 251483 150043 251567
rect 150219 251483 150319 251567
rect 150495 251483 150595 251567
rect 234255 251683 234355 251767
rect 234531 251683 234631 251767
rect 234807 251683 234907 251767
rect 235083 251683 235183 251767
rect 235359 251683 235459 251767
rect 235635 251683 235735 251767
rect 235911 251683 236011 251767
rect 236187 251683 236287 251767
rect 236463 251683 236563 251767
rect 236739 251683 236839 251767
rect 237015 251683 237115 251767
rect 237291 251683 237391 251767
rect 237567 251683 237667 251767
rect 237843 251683 237943 251767
rect 238119 251683 238219 251767
rect 238395 251683 238495 251767
rect 238671 251683 238771 251767
rect 238947 251683 239047 251767
rect 239223 251683 239323 251767
rect 239499 251683 239599 251767
rect 239775 251683 239875 251767
rect 240051 251683 240151 251767
rect 240327 251683 240427 251767
rect 240603 251683 240703 251767
rect 240879 251683 240979 251767
rect 241155 251683 241255 251767
rect 241431 251683 241531 251767
rect 241707 251683 241807 251767
rect 241983 251683 242083 251767
rect 242259 251683 242359 251767
rect 242535 251683 242635 251767
rect 242811 251683 242911 251767
rect 243087 251683 243187 251767
rect 243363 251683 243463 251767
rect 243639 251683 243739 251767
rect 243915 251683 244015 251767
rect 244191 251683 244291 251767
rect 244467 251683 244567 251767
rect 244743 251683 244843 251767
rect 245019 251683 245119 251767
rect 245295 251683 245395 251767
rect 245571 251683 245671 251767
rect 245847 251683 245947 251767
rect 246123 251683 246223 251767
rect 246399 251683 246499 251767
rect 246675 251683 246775 251767
rect 246951 251683 247051 251767
rect 247227 251683 247327 251767
rect 247503 251683 247603 251767
rect 247779 251683 247879 251767
rect 248055 251683 248155 251767
rect 413337 251397 413437 251481
rect 413613 251397 413713 251481
rect 413889 251397 413989 251481
rect 414165 251397 414265 251481
rect 414441 251397 414541 251481
rect 414717 251397 414817 251481
rect 414993 251397 415093 251481
rect 415269 251397 415369 251481
rect 415545 251397 415645 251481
rect 415821 251397 415921 251481
rect 416097 251397 416197 251481
rect 416373 251397 416473 251481
rect 416649 251397 416749 251481
rect 416925 251397 417025 251481
rect 417201 251397 417301 251481
rect 417477 251397 417577 251481
rect 417753 251397 417853 251481
rect 418029 251397 418129 251481
rect 418305 251397 418405 251481
rect 418581 251397 418681 251481
rect 418857 251397 418957 251481
rect 419133 251397 419233 251481
rect 419409 251397 419509 251481
rect 419685 251397 419785 251481
rect 419961 251397 420061 251481
rect 420237 251397 420337 251481
rect 420513 251397 420613 251481
rect 420789 251397 420889 251481
rect 421065 251397 421165 251481
rect 421341 251397 421441 251481
rect 421617 251397 421717 251481
rect 421893 251397 421993 251481
rect 422169 251397 422269 251481
rect 422445 251397 422545 251481
rect 422721 251397 422821 251481
rect 422997 251397 423097 251481
rect 423273 251397 423373 251481
rect 423549 251397 423649 251481
rect 423825 251397 423925 251481
rect 424101 251397 424201 251481
rect 424377 251397 424477 251481
rect 424653 251397 424753 251481
rect 424929 251397 425029 251481
rect 425205 251397 425305 251481
rect 425481 251397 425581 251481
rect 425757 251397 425857 251481
rect 426033 251397 426133 251481
rect 426309 251397 426409 251481
rect 426585 251397 426685 251481
rect 426861 251397 426961 251481
rect 427137 251397 427237 251481
rect 503337 251397 503437 251481
rect 503613 251397 503713 251481
rect 503889 251397 503989 251481
rect 504165 251397 504265 251481
rect 504441 251397 504541 251481
rect 504717 251397 504817 251481
rect 504993 251397 505093 251481
rect 505269 251397 505369 251481
rect 505545 251397 505645 251481
rect 505821 251397 505921 251481
rect 506097 251397 506197 251481
rect 506373 251397 506473 251481
rect 506649 251397 506749 251481
rect 506925 251397 507025 251481
rect 507201 251397 507301 251481
rect 507477 251397 507577 251481
rect 507753 251397 507853 251481
rect 508029 251397 508129 251481
rect 508305 251397 508405 251481
rect 508581 251397 508681 251481
rect 508857 251397 508957 251481
rect 509133 251397 509233 251481
rect 509409 251397 509509 251481
rect 509685 251397 509785 251481
rect 509961 251397 510061 251481
rect 510237 251397 510337 251481
rect 510513 251397 510613 251481
rect 510789 251397 510889 251481
rect 511065 251397 511165 251481
rect 511341 251397 511441 251481
rect 511617 251397 511717 251481
rect 511893 251397 511993 251481
rect 512169 251397 512269 251481
rect 512445 251397 512545 251481
rect 512721 251397 512821 251481
rect 512997 251397 513097 251481
rect 513273 251397 513373 251481
rect 513549 251397 513649 251481
rect 513825 251397 513925 251481
rect 514101 251397 514201 251481
rect 514377 251397 514477 251481
rect 514653 251397 514753 251481
rect 514929 251397 515029 251481
rect 515205 251397 515305 251481
rect 515481 251397 515581 251481
rect 515757 251397 515857 251481
rect 516033 251397 516133 251481
rect 516309 251397 516409 251481
rect 516585 251397 516685 251481
rect 516861 251397 516961 251481
rect 517137 251397 517237 251481
rect 322694 250801 322794 250885
rect 322970 250801 323070 250885
rect 323246 250801 323346 250885
rect 323522 250801 323622 250885
rect 323798 250801 323898 250885
rect 324074 250801 324174 250885
rect 324350 250801 324450 250885
rect 324626 250801 324726 250885
rect 324902 250801 325002 250885
rect 325178 250801 325278 250885
rect 325454 250801 325554 250885
rect 325730 250801 325830 250885
rect 326006 250801 326106 250885
rect 326282 250801 326382 250885
rect 326558 250801 326658 250885
rect 326834 250801 326934 250885
rect 327110 250801 327210 250885
rect 327386 250801 327486 250885
rect 327662 250801 327762 250885
rect 327938 250801 328038 250885
rect 328214 250801 328314 250885
rect 328490 250801 328590 250885
rect 328766 250801 328866 250885
rect 329042 250801 329142 250885
rect 329318 250801 329418 250885
rect 329594 250801 329694 250885
rect 329870 250801 329970 250885
rect 330146 250801 330246 250885
rect 330422 250801 330522 250885
rect 330698 250801 330798 250885
rect 330974 250801 331074 250885
rect 331250 250801 331350 250885
rect 331526 250801 331626 250885
rect 331802 250801 331902 250885
rect 332078 250801 332178 250885
rect 332354 250801 332454 250885
rect 332630 250801 332730 250885
rect 332906 250801 333006 250885
rect 333182 250801 333282 250885
rect 333458 250801 333558 250885
rect 333734 250801 333834 250885
rect 334010 250801 334110 250885
rect 334286 250801 334386 250885
rect 334562 250801 334662 250885
rect 334838 250801 334938 250885
rect 335114 250801 335214 250885
rect 335390 250801 335490 250885
rect 335666 250801 335766 250885
rect 335942 250801 336042 250885
rect 336218 250801 336318 250885
rect 336494 250801 336594 250885
rect 149611 55783 149711 55983
rect 419611 55783 419711 55983
<< mvnmos >>
rect 509423 582417 509523 582617
rect 149621 580493 149721 580693
rect 239621 55493 239721 55693
rect 509621 55493 509721 55693
<< mvpmos >>
rect 419323 657266 419423 657466
rect 329521 580342 329621 580542
rect 149521 145342 149621 145542
rect 419521 145342 419621 145542
<< ndiff >>
rect 329102 657896 329160 657908
rect 329102 657720 329114 657896
rect 329148 657720 329160 657896
rect 329102 657708 329160 657720
rect 329190 657896 329248 657908
rect 329190 657720 329202 657896
rect 329236 657720 329248 657896
rect 329190 657708 329248 657720
rect 509102 657896 509160 657908
rect 509102 657720 509114 657896
rect 509148 657720 509160 657896
rect 509102 657708 509160 657720
rect 509190 657896 509248 657908
rect 509190 657720 509202 657896
rect 509236 657720 509248 657896
rect 509190 657708 509248 657720
rect 149300 655972 149358 655984
rect 149300 655796 149312 655972
rect 149346 655796 149358 655972
rect 149300 655784 149358 655796
rect 149388 655972 149446 655984
rect 149388 655796 149400 655972
rect 149434 655796 149446 655972
rect 149388 655784 149446 655796
rect 239300 580972 239358 580984
rect 239300 580796 239312 580972
rect 239346 580796 239358 580972
rect 239300 580784 239358 580796
rect 239388 580972 239446 580984
rect 239388 580796 239400 580972
rect 239434 580796 239446 580972
rect 239388 580784 239446 580796
rect 239300 145972 239358 145984
rect 239300 145796 239312 145972
rect 239346 145796 239358 145972
rect 239300 145784 239358 145796
rect 239388 145972 239446 145984
rect 239388 145796 239400 145972
rect 239434 145796 239446 145972
rect 239388 145784 239446 145796
rect 509300 145972 509358 145984
rect 509300 145796 509312 145972
rect 509346 145796 509358 145972
rect 509300 145784 509358 145796
rect 509388 145972 509446 145984
rect 509388 145796 509400 145972
rect 509434 145796 509446 145972
rect 509388 145784 509446 145796
rect 59300 55972 59358 55984
rect 59300 55796 59312 55972
rect 59346 55796 59358 55972
rect 59300 55784 59358 55796
rect 59388 55972 59446 55984
rect 59388 55796 59400 55972
rect 59434 55796 59446 55972
rect 59388 55784 59446 55796
rect 329300 55972 329358 55984
rect 329300 55796 329312 55972
rect 329346 55796 329358 55972
rect 329300 55784 329358 55796
rect 329388 55972 329446 55984
rect 329388 55796 329400 55972
rect 329434 55796 329446 55972
rect 329388 55784 329446 55796
<< pdiff >>
rect 239283 655934 239341 655946
rect 239283 655758 239295 655934
rect 239329 655758 239341 655934
rect 239283 655746 239341 655758
rect 239371 655934 239429 655946
rect 239371 655758 239383 655934
rect 239417 655758 239429 655934
rect 239371 655746 239429 655758
rect 59283 145934 59341 145946
rect 59283 145758 59295 145934
rect 59329 145758 59341 145934
rect 59283 145746 59341 145758
rect 59371 145934 59429 145946
rect 59371 145758 59383 145934
rect 59417 145758 59429 145934
rect 59371 145746 59429 145758
rect 329283 145934 329341 145946
rect 329283 145758 329295 145934
rect 329329 145758 329341 145934
rect 329283 145746 329341 145758
rect 329371 145934 329429 145946
rect 329371 145758 329383 145934
rect 329417 145758 329429 145934
rect 329371 145746 329429 145758
<< mvndiff >>
rect 59553 655971 59611 655983
rect 59553 655795 59565 655971
rect 59599 655795 59611 655971
rect 59553 655783 59611 655795
rect 59711 655971 59769 655983
rect 59711 655795 59723 655971
rect 59757 655795 59769 655971
rect 59711 655783 59769 655795
rect 419355 582895 419413 582907
rect 419355 582719 419367 582895
rect 419401 582719 419413 582895
rect 419355 582707 419413 582719
rect 419513 582895 419571 582907
rect 419513 582719 419525 582895
rect 419559 582719 419571 582895
rect 419513 582707 419571 582719
rect 509365 582605 509423 582617
rect 509365 582429 509377 582605
rect 509411 582429 509423 582605
rect 509365 582417 509423 582429
rect 509523 582605 509581 582617
rect 509523 582429 509535 582605
rect 509569 582429 509581 582605
rect 509523 582417 509581 582429
rect 59553 580971 59611 580983
rect 59553 580795 59565 580971
rect 59599 580795 59611 580971
rect 59553 580783 59611 580795
rect 59711 580971 59769 580983
rect 59711 580795 59723 580971
rect 59757 580795 59769 580971
rect 59711 580783 59769 580795
rect 149563 580681 149621 580693
rect 149563 580505 149575 580681
rect 149609 580505 149621 580681
rect 149563 580493 149621 580505
rect 149721 580681 149779 580693
rect 149721 580505 149733 580681
rect 149767 580505 149779 580681
rect 149721 580493 149779 580505
rect 58829 491759 58887 491771
rect 58829 491699 58841 491759
rect 58875 491699 58887 491759
rect 58829 491687 58887 491699
rect 58987 491759 59045 491771
rect 58987 491699 58999 491759
rect 59033 491699 59045 491759
rect 58987 491687 59045 491699
rect 59105 491759 59163 491771
rect 59105 491699 59117 491759
rect 59151 491699 59163 491759
rect 59105 491687 59163 491699
rect 59263 491759 59321 491771
rect 59263 491699 59275 491759
rect 59309 491699 59321 491759
rect 59263 491687 59321 491699
rect 59381 491759 59439 491771
rect 59381 491699 59393 491759
rect 59427 491699 59439 491759
rect 59381 491687 59439 491699
rect 59539 491759 59597 491771
rect 59539 491699 59551 491759
rect 59585 491699 59597 491759
rect 59539 491687 59597 491699
rect 59657 491759 59715 491771
rect 59657 491699 59669 491759
rect 59703 491699 59715 491759
rect 59657 491687 59715 491699
rect 59815 491759 59873 491771
rect 59815 491699 59827 491759
rect 59861 491699 59873 491759
rect 59815 491687 59873 491699
rect 59933 491759 59991 491771
rect 59933 491699 59945 491759
rect 59979 491699 59991 491759
rect 59933 491687 59991 491699
rect 60091 491759 60149 491771
rect 60091 491699 60103 491759
rect 60137 491699 60149 491759
rect 60091 491687 60149 491699
rect 60209 491759 60267 491771
rect 60209 491699 60221 491759
rect 60255 491699 60267 491759
rect 60209 491687 60267 491699
rect 60367 491759 60425 491771
rect 60367 491699 60379 491759
rect 60413 491699 60425 491759
rect 60367 491687 60425 491699
rect 60485 491759 60543 491771
rect 60485 491699 60497 491759
rect 60531 491699 60543 491759
rect 60485 491687 60543 491699
rect 60643 491759 60701 491771
rect 60643 491699 60655 491759
rect 60689 491699 60701 491759
rect 60643 491687 60701 491699
rect 60761 491759 60819 491771
rect 60761 491699 60773 491759
rect 60807 491699 60819 491759
rect 60761 491687 60819 491699
rect 60919 491759 60977 491771
rect 60919 491699 60931 491759
rect 60965 491699 60977 491759
rect 60919 491687 60977 491699
rect 61037 491759 61095 491771
rect 61037 491699 61049 491759
rect 61083 491699 61095 491759
rect 61037 491687 61095 491699
rect 61195 491759 61253 491771
rect 61195 491699 61207 491759
rect 61241 491699 61253 491759
rect 61195 491687 61253 491699
rect 61313 491759 61371 491771
rect 61313 491699 61325 491759
rect 61359 491699 61371 491759
rect 61313 491687 61371 491699
rect 61471 491759 61529 491771
rect 61471 491699 61483 491759
rect 61517 491699 61529 491759
rect 61471 491687 61529 491699
rect 323819 492147 323877 492159
rect 323819 492087 323831 492147
rect 323865 492087 323877 492147
rect 323819 492075 323877 492087
rect 323977 492147 324035 492159
rect 323977 492087 323989 492147
rect 324023 492087 324035 492147
rect 323977 492075 324035 492087
rect 324095 492147 324153 492159
rect 324095 492087 324107 492147
rect 324141 492087 324153 492147
rect 324095 492075 324153 492087
rect 324253 492147 324311 492159
rect 324253 492087 324265 492147
rect 324299 492087 324311 492147
rect 324253 492075 324311 492087
rect 324371 492147 324429 492159
rect 324371 492087 324383 492147
rect 324417 492087 324429 492147
rect 324371 492075 324429 492087
rect 324529 492147 324587 492159
rect 324529 492087 324541 492147
rect 324575 492087 324587 492147
rect 324529 492075 324587 492087
rect 324647 492147 324705 492159
rect 324647 492087 324659 492147
rect 324693 492087 324705 492147
rect 324647 492075 324705 492087
rect 324805 492147 324863 492159
rect 324805 492087 324817 492147
rect 324851 492087 324863 492147
rect 324805 492075 324863 492087
rect 324923 492147 324981 492159
rect 324923 492087 324935 492147
rect 324969 492087 324981 492147
rect 324923 492075 324981 492087
rect 325081 492147 325139 492159
rect 325081 492087 325093 492147
rect 325127 492087 325139 492147
rect 325081 492075 325139 492087
rect 325199 492147 325257 492159
rect 325199 492087 325211 492147
rect 325245 492087 325257 492147
rect 325199 492075 325257 492087
rect 325357 492147 325415 492159
rect 325357 492087 325369 492147
rect 325403 492087 325415 492147
rect 325357 492075 325415 492087
rect 325475 492147 325533 492159
rect 325475 492087 325487 492147
rect 325521 492087 325533 492147
rect 325475 492075 325533 492087
rect 325633 492147 325691 492159
rect 325633 492087 325645 492147
rect 325679 492087 325691 492147
rect 325633 492075 325691 492087
rect 325751 492147 325809 492159
rect 325751 492087 325763 492147
rect 325797 492087 325809 492147
rect 325751 492075 325809 492087
rect 325909 492147 325967 492159
rect 325909 492087 325921 492147
rect 325955 492087 325967 492147
rect 325909 492075 325967 492087
rect 326027 492147 326085 492159
rect 326027 492087 326039 492147
rect 326073 492087 326085 492147
rect 326027 492075 326085 492087
rect 326185 492147 326243 492159
rect 326185 492087 326197 492147
rect 326231 492087 326243 492147
rect 326185 492075 326243 492087
rect 326303 492147 326361 492159
rect 326303 492087 326315 492147
rect 326349 492087 326361 492147
rect 326303 492075 326361 492087
rect 326461 492147 326519 492159
rect 326461 492087 326473 492147
rect 326507 492087 326519 492147
rect 326461 492075 326519 492087
rect 326579 492147 326637 492159
rect 326579 492087 326591 492147
rect 326625 492087 326637 492147
rect 326579 492075 326637 492087
rect 326737 492147 326795 492159
rect 326737 492087 326749 492147
rect 326783 492087 326795 492147
rect 326737 492075 326795 492087
rect 326855 492147 326913 492159
rect 326855 492087 326867 492147
rect 326901 492087 326913 492147
rect 326855 492075 326913 492087
rect 327013 492147 327071 492159
rect 327013 492087 327025 492147
rect 327059 492087 327071 492147
rect 327013 492075 327071 492087
rect 327131 492147 327189 492159
rect 327131 492087 327143 492147
rect 327177 492087 327189 492147
rect 327131 492075 327189 492087
rect 327289 492147 327347 492159
rect 327289 492087 327301 492147
rect 327335 492087 327347 492147
rect 327289 492075 327347 492087
rect 327407 492147 327465 492159
rect 327407 492087 327419 492147
rect 327453 492087 327465 492147
rect 327407 492075 327465 492087
rect 327565 492147 327623 492159
rect 327565 492087 327577 492147
rect 327611 492087 327623 492147
rect 327565 492075 327623 492087
rect 327683 492147 327741 492159
rect 327683 492087 327695 492147
rect 327729 492087 327741 492147
rect 327683 492075 327741 492087
rect 327841 492147 327899 492159
rect 327841 492087 327853 492147
rect 327887 492087 327899 492147
rect 327841 492075 327899 492087
rect 327959 492147 328017 492159
rect 327959 492087 327971 492147
rect 328005 492087 328017 492147
rect 327959 492075 328017 492087
rect 328117 492147 328175 492159
rect 328117 492087 328129 492147
rect 328163 492087 328175 492147
rect 328117 492075 328175 492087
rect 328235 492147 328293 492159
rect 328235 492087 328247 492147
rect 328281 492087 328293 492147
rect 328235 492075 328293 492087
rect 328393 492147 328451 492159
rect 328393 492087 328405 492147
rect 328439 492087 328451 492147
rect 328393 492075 328451 492087
rect 328511 492147 328569 492159
rect 328511 492087 328523 492147
rect 328557 492087 328569 492147
rect 328511 492075 328569 492087
rect 328669 492147 328727 492159
rect 328669 492087 328681 492147
rect 328715 492087 328727 492147
rect 328669 492075 328727 492087
rect 328787 492147 328845 492159
rect 328787 492087 328799 492147
rect 328833 492087 328845 492147
rect 328787 492075 328845 492087
rect 328945 492147 329003 492159
rect 328945 492087 328957 492147
rect 328991 492087 329003 492147
rect 328945 492075 329003 492087
rect 329063 492147 329121 492159
rect 329063 492087 329075 492147
rect 329109 492087 329121 492147
rect 329063 492075 329121 492087
rect 329221 492147 329279 492159
rect 329221 492087 329233 492147
rect 329267 492087 329279 492147
rect 329221 492075 329279 492087
rect 329339 492147 329397 492159
rect 329339 492087 329351 492147
rect 329385 492087 329397 492147
rect 329339 492075 329397 492087
rect 329497 492147 329555 492159
rect 329497 492087 329509 492147
rect 329543 492087 329555 492147
rect 329497 492075 329555 492087
rect 329615 492147 329673 492159
rect 329615 492087 329627 492147
rect 329661 492087 329673 492147
rect 329615 492075 329673 492087
rect 329773 492147 329831 492159
rect 329773 492087 329785 492147
rect 329819 492087 329831 492147
rect 329773 492075 329831 492087
rect 329891 492147 329949 492159
rect 329891 492087 329903 492147
rect 329937 492087 329949 492147
rect 329891 492075 329949 492087
rect 330049 492147 330107 492159
rect 330049 492087 330061 492147
rect 330095 492087 330107 492147
rect 330049 492075 330107 492087
rect 330167 492147 330225 492159
rect 330167 492087 330179 492147
rect 330213 492087 330225 492147
rect 330167 492075 330225 492087
rect 330325 492147 330383 492159
rect 330325 492087 330337 492147
rect 330371 492087 330383 492147
rect 330325 492075 330383 492087
rect 330443 492147 330501 492159
rect 330443 492087 330455 492147
rect 330489 492087 330501 492147
rect 330443 492075 330501 492087
rect 330601 492147 330659 492159
rect 330601 492087 330613 492147
rect 330647 492087 330659 492147
rect 330601 492075 330659 492087
rect 330719 492147 330777 492159
rect 330719 492087 330731 492147
rect 330765 492087 330777 492147
rect 330719 492075 330777 492087
rect 330877 492147 330935 492159
rect 330877 492087 330889 492147
rect 330923 492087 330935 492147
rect 330877 492075 330935 492087
rect 330995 492147 331053 492159
rect 330995 492087 331007 492147
rect 331041 492087 331053 492147
rect 330995 492075 331053 492087
rect 331153 492147 331211 492159
rect 331153 492087 331165 492147
rect 331199 492087 331211 492147
rect 331153 492075 331211 492087
rect 331271 492147 331329 492159
rect 331271 492087 331283 492147
rect 331317 492087 331329 492147
rect 331271 492075 331329 492087
rect 331429 492147 331487 492159
rect 331429 492087 331441 492147
rect 331475 492087 331487 492147
rect 331429 492075 331487 492087
rect 331547 492147 331605 492159
rect 331547 492087 331559 492147
rect 331593 492087 331605 492147
rect 331547 492075 331605 492087
rect 331705 492147 331763 492159
rect 331705 492087 331717 492147
rect 331751 492087 331763 492147
rect 331705 492075 331763 492087
rect 331823 492147 331881 492159
rect 331823 492087 331835 492147
rect 331869 492087 331881 492147
rect 331823 492075 331881 492087
rect 331981 492147 332039 492159
rect 331981 492087 331993 492147
rect 332027 492087 332039 492147
rect 331981 492075 332039 492087
rect 332099 492147 332157 492159
rect 332099 492087 332111 492147
rect 332145 492087 332157 492147
rect 332099 492075 332157 492087
rect 332257 492147 332315 492159
rect 332257 492087 332269 492147
rect 332303 492087 332315 492147
rect 332257 492075 332315 492087
rect 332375 492147 332433 492159
rect 332375 492087 332387 492147
rect 332421 492087 332433 492147
rect 332375 492075 332433 492087
rect 332533 492147 332591 492159
rect 332533 492087 332545 492147
rect 332579 492087 332591 492147
rect 332533 492075 332591 492087
rect 332651 492147 332709 492159
rect 332651 492087 332663 492147
rect 332697 492087 332709 492147
rect 332651 492075 332709 492087
rect 332809 492147 332867 492159
rect 332809 492087 332821 492147
rect 332855 492087 332867 492147
rect 332809 492075 332867 492087
rect 332927 492147 332985 492159
rect 332927 492087 332939 492147
rect 332973 492087 332985 492147
rect 332927 492075 332985 492087
rect 333085 492147 333143 492159
rect 333085 492087 333097 492147
rect 333131 492087 333143 492147
rect 333085 492075 333143 492087
rect 333203 492147 333261 492159
rect 333203 492087 333215 492147
rect 333249 492087 333261 492147
rect 333203 492075 333261 492087
rect 333361 492147 333419 492159
rect 333361 492087 333373 492147
rect 333407 492087 333419 492147
rect 333361 492075 333419 492087
rect 333479 492147 333537 492159
rect 333479 492087 333491 492147
rect 333525 492087 333537 492147
rect 333479 492075 333537 492087
rect 333637 492147 333695 492159
rect 333637 492087 333649 492147
rect 333683 492087 333695 492147
rect 333637 492075 333695 492087
rect 333755 492147 333813 492159
rect 333755 492087 333767 492147
rect 333801 492087 333813 492147
rect 333755 492075 333813 492087
rect 333913 492147 333971 492159
rect 333913 492087 333925 492147
rect 333959 492087 333971 492147
rect 333913 492075 333971 492087
rect 334031 492147 334089 492159
rect 334031 492087 334043 492147
rect 334077 492087 334089 492147
rect 334031 492075 334089 492087
rect 334189 492147 334247 492159
rect 334189 492087 334201 492147
rect 334235 492087 334247 492147
rect 334189 492075 334247 492087
rect 334307 492147 334365 492159
rect 334307 492087 334319 492147
rect 334353 492087 334365 492147
rect 334307 492075 334365 492087
rect 334465 492147 334523 492159
rect 334465 492087 334477 492147
rect 334511 492087 334523 492147
rect 334465 492075 334523 492087
rect 334583 492147 334641 492159
rect 334583 492087 334595 492147
rect 334629 492087 334641 492147
rect 334583 492075 334641 492087
rect 334741 492147 334799 492159
rect 334741 492087 334753 492147
rect 334787 492087 334799 492147
rect 334741 492075 334799 492087
rect 334859 492147 334917 492159
rect 334859 492087 334871 492147
rect 334905 492087 334917 492147
rect 334859 492075 334917 492087
rect 335017 492147 335075 492159
rect 335017 492087 335029 492147
rect 335063 492087 335075 492147
rect 335017 492075 335075 492087
rect 335135 492147 335193 492159
rect 335135 492087 335147 492147
rect 335181 492087 335193 492147
rect 335135 492075 335193 492087
rect 335293 492147 335351 492159
rect 335293 492087 335305 492147
rect 335339 492087 335351 492147
rect 335293 492075 335351 492087
rect 335411 492147 335469 492159
rect 335411 492087 335423 492147
rect 335457 492087 335469 492147
rect 335411 492075 335469 492087
rect 335569 492147 335627 492159
rect 335569 492087 335581 492147
rect 335615 492087 335627 492147
rect 335569 492075 335627 492087
rect 335687 492147 335745 492159
rect 335687 492087 335699 492147
rect 335733 492087 335745 492147
rect 335687 492075 335745 492087
rect 335845 492147 335903 492159
rect 335845 492087 335857 492147
rect 335891 492087 335903 492147
rect 335845 492075 335903 492087
rect 335963 492147 336021 492159
rect 335963 492087 335975 492147
rect 336009 492087 336021 492147
rect 335963 492075 336021 492087
rect 336121 492147 336179 492159
rect 336121 492087 336133 492147
rect 336167 492087 336179 492147
rect 336121 492075 336179 492087
rect 336239 492147 336297 492159
rect 336239 492087 336251 492147
rect 336285 492087 336297 492147
rect 336239 492075 336297 492087
rect 336397 492147 336455 492159
rect 336397 492087 336409 492147
rect 336443 492087 336455 492147
rect 336397 492075 336455 492087
rect 336515 492147 336573 492159
rect 336515 492087 336527 492147
rect 336561 492087 336573 492147
rect 336515 492075 336573 492087
rect 336673 492147 336731 492159
rect 336673 492087 336685 492147
rect 336719 492087 336731 492147
rect 336673 492075 336731 492087
rect 336791 492147 336849 492159
rect 336791 492087 336803 492147
rect 336837 492087 336849 492147
rect 336791 492075 336849 492087
rect 336949 492147 337007 492159
rect 336949 492087 336961 492147
rect 336995 492087 337007 492147
rect 336949 492075 337007 492087
rect 337067 492147 337125 492159
rect 337067 492087 337079 492147
rect 337113 492087 337125 492147
rect 337067 492075 337125 492087
rect 337225 492147 337283 492159
rect 337225 492087 337237 492147
rect 337271 492087 337283 492147
rect 337225 492075 337283 492087
rect 337343 492147 337401 492159
rect 337343 492087 337355 492147
rect 337389 492087 337401 492147
rect 337343 492075 337401 492087
rect 337501 492147 337559 492159
rect 337501 492087 337513 492147
rect 337547 492087 337559 492147
rect 337501 492075 337559 492087
rect 337619 492147 337677 492159
rect 337619 492087 337631 492147
rect 337665 492087 337677 492147
rect 337619 492075 337677 492087
rect 337777 492147 337835 492159
rect 337777 492087 337789 492147
rect 337823 492087 337835 492147
rect 337777 492075 337835 492087
rect 143279 491469 143337 491481
rect 143279 491409 143291 491469
rect 143325 491409 143337 491469
rect 143279 491397 143337 491409
rect 143437 491469 143495 491481
rect 143437 491409 143449 491469
rect 143483 491409 143495 491469
rect 143437 491397 143495 491409
rect 143555 491469 143613 491481
rect 143555 491409 143567 491469
rect 143601 491409 143613 491469
rect 143555 491397 143613 491409
rect 143713 491469 143771 491481
rect 143713 491409 143725 491469
rect 143759 491409 143771 491469
rect 143713 491397 143771 491409
rect 143831 491469 143889 491481
rect 143831 491409 143843 491469
rect 143877 491409 143889 491469
rect 143831 491397 143889 491409
rect 143989 491469 144047 491481
rect 143989 491409 144001 491469
rect 144035 491409 144047 491469
rect 143989 491397 144047 491409
rect 144107 491469 144165 491481
rect 144107 491409 144119 491469
rect 144153 491409 144165 491469
rect 144107 491397 144165 491409
rect 144265 491469 144323 491481
rect 144265 491409 144277 491469
rect 144311 491409 144323 491469
rect 144265 491397 144323 491409
rect 144383 491469 144441 491481
rect 144383 491409 144395 491469
rect 144429 491409 144441 491469
rect 144383 491397 144441 491409
rect 144541 491469 144599 491481
rect 144541 491409 144553 491469
rect 144587 491409 144599 491469
rect 144541 491397 144599 491409
rect 144659 491469 144717 491481
rect 144659 491409 144671 491469
rect 144705 491409 144717 491469
rect 144659 491397 144717 491409
rect 144817 491469 144875 491481
rect 144817 491409 144829 491469
rect 144863 491409 144875 491469
rect 144817 491397 144875 491409
rect 144935 491469 144993 491481
rect 144935 491409 144947 491469
rect 144981 491409 144993 491469
rect 144935 491397 144993 491409
rect 145093 491469 145151 491481
rect 145093 491409 145105 491469
rect 145139 491409 145151 491469
rect 145093 491397 145151 491409
rect 145211 491469 145269 491481
rect 145211 491409 145223 491469
rect 145257 491409 145269 491469
rect 145211 491397 145269 491409
rect 145369 491469 145427 491481
rect 145369 491409 145381 491469
rect 145415 491409 145427 491469
rect 145369 491397 145427 491409
rect 145487 491469 145545 491481
rect 145487 491409 145499 491469
rect 145533 491409 145545 491469
rect 145487 491397 145545 491409
rect 145645 491469 145703 491481
rect 145645 491409 145657 491469
rect 145691 491409 145703 491469
rect 145645 491397 145703 491409
rect 145763 491469 145821 491481
rect 145763 491409 145775 491469
rect 145809 491409 145821 491469
rect 145763 491397 145821 491409
rect 145921 491469 145979 491481
rect 145921 491409 145933 491469
rect 145967 491409 145979 491469
rect 145921 491397 145979 491409
rect 146039 491469 146097 491481
rect 146039 491409 146051 491469
rect 146085 491409 146097 491469
rect 146039 491397 146097 491409
rect 146197 491469 146255 491481
rect 146197 491409 146209 491469
rect 146243 491409 146255 491469
rect 146197 491397 146255 491409
rect 146315 491469 146373 491481
rect 146315 491409 146327 491469
rect 146361 491409 146373 491469
rect 146315 491397 146373 491409
rect 146473 491469 146531 491481
rect 146473 491409 146485 491469
rect 146519 491409 146531 491469
rect 146473 491397 146531 491409
rect 146591 491469 146649 491481
rect 146591 491409 146603 491469
rect 146637 491409 146649 491469
rect 146591 491397 146649 491409
rect 146749 491469 146807 491481
rect 146749 491409 146761 491469
rect 146795 491409 146807 491469
rect 146749 491397 146807 491409
rect 146867 491469 146925 491481
rect 146867 491409 146879 491469
rect 146913 491409 146925 491469
rect 146867 491397 146925 491409
rect 147025 491469 147083 491481
rect 147025 491409 147037 491469
rect 147071 491409 147083 491469
rect 147025 491397 147083 491409
rect 147143 491469 147201 491481
rect 147143 491409 147155 491469
rect 147189 491409 147201 491469
rect 147143 491397 147201 491409
rect 147301 491469 147359 491481
rect 147301 491409 147313 491469
rect 147347 491409 147359 491469
rect 147301 491397 147359 491409
rect 147419 491469 147477 491481
rect 147419 491409 147431 491469
rect 147465 491409 147477 491469
rect 147419 491397 147477 491409
rect 147577 491469 147635 491481
rect 147577 491409 147589 491469
rect 147623 491409 147635 491469
rect 147577 491397 147635 491409
rect 147695 491469 147753 491481
rect 147695 491409 147707 491469
rect 147741 491409 147753 491469
rect 147695 491397 147753 491409
rect 147853 491469 147911 491481
rect 147853 491409 147865 491469
rect 147899 491409 147911 491469
rect 147853 491397 147911 491409
rect 147971 491469 148029 491481
rect 147971 491409 147983 491469
rect 148017 491409 148029 491469
rect 147971 491397 148029 491409
rect 148129 491469 148187 491481
rect 148129 491409 148141 491469
rect 148175 491409 148187 491469
rect 148129 491397 148187 491409
rect 148247 491469 148305 491481
rect 148247 491409 148259 491469
rect 148293 491409 148305 491469
rect 148247 491397 148305 491409
rect 148405 491469 148463 491481
rect 148405 491409 148417 491469
rect 148451 491409 148463 491469
rect 148405 491397 148463 491409
rect 148523 491469 148581 491481
rect 148523 491409 148535 491469
rect 148569 491409 148581 491469
rect 148523 491397 148581 491409
rect 148681 491469 148739 491481
rect 148681 491409 148693 491469
rect 148727 491409 148739 491469
rect 148681 491397 148739 491409
rect 148799 491469 148857 491481
rect 148799 491409 148811 491469
rect 148845 491409 148857 491469
rect 148799 491397 148857 491409
rect 148957 491469 149015 491481
rect 148957 491409 148969 491469
rect 149003 491409 149015 491469
rect 148957 491397 149015 491409
rect 149075 491469 149133 491481
rect 149075 491409 149087 491469
rect 149121 491409 149133 491469
rect 149075 491397 149133 491409
rect 149233 491469 149291 491481
rect 149233 491409 149245 491469
rect 149279 491409 149291 491469
rect 149233 491397 149291 491409
rect 149351 491469 149409 491481
rect 149351 491409 149363 491469
rect 149397 491409 149409 491469
rect 149351 491397 149409 491409
rect 149509 491469 149567 491481
rect 149509 491409 149521 491469
rect 149555 491409 149567 491469
rect 149509 491397 149567 491409
rect 149627 491469 149685 491481
rect 149627 491409 149639 491469
rect 149673 491409 149685 491469
rect 149627 491397 149685 491409
rect 149785 491469 149843 491481
rect 149785 491409 149797 491469
rect 149831 491409 149843 491469
rect 149785 491397 149843 491409
rect 149903 491469 149961 491481
rect 149903 491409 149915 491469
rect 149949 491409 149961 491469
rect 149903 491397 149961 491409
rect 150061 491469 150119 491481
rect 150061 491409 150073 491469
rect 150107 491409 150119 491469
rect 150061 491397 150119 491409
rect 150179 491469 150237 491481
rect 150179 491409 150191 491469
rect 150225 491409 150237 491469
rect 150179 491397 150237 491409
rect 150337 491469 150395 491481
rect 150337 491409 150349 491469
rect 150383 491409 150395 491469
rect 150337 491397 150395 491409
rect 150455 491469 150513 491481
rect 150455 491409 150467 491469
rect 150501 491409 150513 491469
rect 150455 491397 150513 491409
rect 150613 491469 150671 491481
rect 150613 491409 150625 491469
rect 150659 491409 150671 491469
rect 150613 491397 150671 491409
rect 150731 491469 150789 491481
rect 150731 491409 150743 491469
rect 150777 491409 150789 491469
rect 150731 491397 150789 491409
rect 150889 491469 150947 491481
rect 150889 491409 150901 491469
rect 150935 491409 150947 491469
rect 150889 491397 150947 491409
rect 151007 491469 151065 491481
rect 151007 491409 151019 491469
rect 151053 491409 151065 491469
rect 151007 491397 151065 491409
rect 151165 491469 151223 491481
rect 151165 491409 151177 491469
rect 151211 491409 151223 491469
rect 151165 491397 151223 491409
rect 151283 491469 151341 491481
rect 151283 491409 151295 491469
rect 151329 491409 151341 491469
rect 151283 491397 151341 491409
rect 151441 491469 151499 491481
rect 151441 491409 151453 491469
rect 151487 491409 151499 491469
rect 151441 491397 151499 491409
rect 151559 491469 151617 491481
rect 151559 491409 151571 491469
rect 151605 491409 151617 491469
rect 151559 491397 151617 491409
rect 151717 491469 151775 491481
rect 151717 491409 151729 491469
rect 151763 491409 151775 491469
rect 151717 491397 151775 491409
rect 151835 491469 151893 491481
rect 151835 491409 151847 491469
rect 151881 491409 151893 491469
rect 151835 491397 151893 491409
rect 151993 491469 152051 491481
rect 151993 491409 152005 491469
rect 152039 491409 152051 491469
rect 151993 491397 152051 491409
rect 152111 491469 152169 491481
rect 152111 491409 152123 491469
rect 152157 491409 152169 491469
rect 152111 491397 152169 491409
rect 152269 491469 152327 491481
rect 152269 491409 152281 491469
rect 152315 491409 152327 491469
rect 152269 491397 152327 491409
rect 152387 491469 152445 491481
rect 152387 491409 152399 491469
rect 152433 491409 152445 491469
rect 152387 491397 152445 491409
rect 152545 491469 152603 491481
rect 152545 491409 152557 491469
rect 152591 491409 152603 491469
rect 152545 491397 152603 491409
rect 152663 491469 152721 491481
rect 152663 491409 152675 491469
rect 152709 491409 152721 491469
rect 152663 491397 152721 491409
rect 152821 491469 152879 491481
rect 152821 491409 152833 491469
rect 152867 491409 152879 491469
rect 152821 491397 152879 491409
rect 152939 491469 152997 491481
rect 152939 491409 152951 491469
rect 152985 491409 152997 491469
rect 152939 491397 152997 491409
rect 153097 491469 153155 491481
rect 153097 491409 153109 491469
rect 153143 491409 153155 491469
rect 153097 491397 153155 491409
rect 153215 491469 153273 491481
rect 153215 491409 153227 491469
rect 153261 491409 153273 491469
rect 153215 491397 153273 491409
rect 153373 491469 153431 491481
rect 153373 491409 153385 491469
rect 153419 491409 153431 491469
rect 153373 491397 153431 491409
rect 153491 491469 153549 491481
rect 153491 491409 153503 491469
rect 153537 491409 153549 491469
rect 153491 491397 153549 491409
rect 153649 491469 153707 491481
rect 153649 491409 153661 491469
rect 153695 491409 153707 491469
rect 153649 491397 153707 491409
rect 153767 491469 153825 491481
rect 153767 491409 153779 491469
rect 153813 491409 153825 491469
rect 153767 491397 153825 491409
rect 153925 491469 153983 491481
rect 153925 491409 153937 491469
rect 153971 491409 153983 491469
rect 153925 491397 153983 491409
rect 154043 491469 154101 491481
rect 154043 491409 154055 491469
rect 154089 491409 154101 491469
rect 154043 491397 154101 491409
rect 154201 491469 154259 491481
rect 154201 491409 154213 491469
rect 154247 491409 154259 491469
rect 154201 491397 154259 491409
rect 154319 491469 154377 491481
rect 154319 491409 154331 491469
rect 154365 491409 154377 491469
rect 154319 491397 154377 491409
rect 154477 491469 154535 491481
rect 154477 491409 154489 491469
rect 154523 491409 154535 491469
rect 154477 491397 154535 491409
rect 154595 491469 154653 491481
rect 154595 491409 154607 491469
rect 154641 491409 154653 491469
rect 154595 491397 154653 491409
rect 154753 491469 154811 491481
rect 154753 491409 154765 491469
rect 154799 491409 154811 491469
rect 154753 491397 154811 491409
rect 154871 491469 154929 491481
rect 154871 491409 154883 491469
rect 154917 491409 154929 491469
rect 154871 491397 154929 491409
rect 155029 491469 155087 491481
rect 155029 491409 155041 491469
rect 155075 491409 155087 491469
rect 155029 491397 155087 491409
rect 155147 491469 155205 491481
rect 155147 491409 155159 491469
rect 155193 491409 155205 491469
rect 155147 491397 155205 491409
rect 155305 491469 155363 491481
rect 155305 491409 155317 491469
rect 155351 491409 155363 491469
rect 155305 491397 155363 491409
rect 155423 491469 155481 491481
rect 155423 491409 155435 491469
rect 155469 491409 155481 491469
rect 155423 491397 155481 491409
rect 155581 491469 155639 491481
rect 155581 491409 155593 491469
rect 155627 491409 155639 491469
rect 155581 491397 155639 491409
rect 155699 491469 155757 491481
rect 155699 491409 155711 491469
rect 155745 491409 155757 491469
rect 155699 491397 155757 491409
rect 155857 491469 155915 491481
rect 155857 491409 155869 491469
rect 155903 491409 155915 491469
rect 155857 491397 155915 491409
rect 155975 491469 156033 491481
rect 155975 491409 155987 491469
rect 156021 491409 156033 491469
rect 155975 491397 156033 491409
rect 156133 491469 156191 491481
rect 156133 491409 156145 491469
rect 156179 491409 156191 491469
rect 156133 491397 156191 491409
rect 156251 491469 156309 491481
rect 156251 491409 156263 491469
rect 156297 491409 156309 491469
rect 156251 491397 156309 491409
rect 156409 491469 156467 491481
rect 156409 491409 156421 491469
rect 156455 491409 156467 491469
rect 156409 491397 156467 491409
rect 156527 491469 156585 491481
rect 156527 491409 156539 491469
rect 156573 491409 156585 491469
rect 156527 491397 156585 491409
rect 156685 491469 156743 491481
rect 156685 491409 156697 491469
rect 156731 491409 156743 491469
rect 156685 491397 156743 491409
rect 156803 491469 156861 491481
rect 156803 491409 156815 491469
rect 156849 491409 156861 491469
rect 156803 491397 156861 491409
rect 156961 491469 157019 491481
rect 156961 491409 156973 491469
rect 157007 491409 157019 491469
rect 156961 491397 157019 491409
rect 157079 491469 157137 491481
rect 157079 491409 157091 491469
rect 157125 491409 157137 491469
rect 157079 491397 157137 491409
rect 157237 491469 157295 491481
rect 157237 491409 157249 491469
rect 157283 491409 157295 491469
rect 157237 491397 157295 491409
rect 418828 491431 418886 491443
rect 418828 491371 418840 491431
rect 418874 491371 418886 491431
rect 418828 491359 418886 491371
rect 418986 491431 419044 491443
rect 418986 491371 418998 491431
rect 419032 491371 419044 491431
rect 418986 491359 419044 491371
rect 419104 491431 419162 491443
rect 419104 491371 419116 491431
rect 419150 491371 419162 491431
rect 419104 491359 419162 491371
rect 419262 491431 419320 491443
rect 419262 491371 419274 491431
rect 419308 491371 419320 491431
rect 419262 491359 419320 491371
rect 419380 491431 419438 491443
rect 419380 491371 419392 491431
rect 419426 491371 419438 491431
rect 419380 491359 419438 491371
rect 419538 491431 419596 491443
rect 419538 491371 419550 491431
rect 419584 491371 419596 491431
rect 419538 491359 419596 491371
rect 419656 491431 419714 491443
rect 419656 491371 419668 491431
rect 419702 491371 419714 491431
rect 419656 491359 419714 491371
rect 419814 491431 419872 491443
rect 419814 491371 419826 491431
rect 419860 491371 419872 491431
rect 419814 491359 419872 491371
rect 419932 491431 419990 491443
rect 419932 491371 419944 491431
rect 419978 491371 419990 491431
rect 419932 491359 419990 491371
rect 420090 491431 420148 491443
rect 420090 491371 420102 491431
rect 420136 491371 420148 491431
rect 420090 491359 420148 491371
rect 508829 491759 508887 491771
rect 508829 491699 508841 491759
rect 508875 491699 508887 491759
rect 508829 491687 508887 491699
rect 508987 491759 509045 491771
rect 508987 491699 508999 491759
rect 509033 491699 509045 491759
rect 508987 491687 509045 491699
rect 509105 491759 509163 491771
rect 509105 491699 509117 491759
rect 509151 491699 509163 491759
rect 509105 491687 509163 491699
rect 509263 491759 509321 491771
rect 509263 491699 509275 491759
rect 509309 491699 509321 491759
rect 509263 491687 509321 491699
rect 509381 491759 509439 491771
rect 509381 491699 509393 491759
rect 509427 491699 509439 491759
rect 509381 491687 509439 491699
rect 509539 491759 509597 491771
rect 509539 491699 509551 491759
rect 509585 491699 509597 491759
rect 509539 491687 509597 491699
rect 509657 491759 509715 491771
rect 509657 491699 509669 491759
rect 509703 491699 509715 491759
rect 509657 491687 509715 491699
rect 509815 491759 509873 491771
rect 509815 491699 509827 491759
rect 509861 491699 509873 491759
rect 509815 491687 509873 491699
rect 509933 491759 509991 491771
rect 509933 491699 509945 491759
rect 509979 491699 509991 491759
rect 509933 491687 509991 491699
rect 510091 491759 510149 491771
rect 510091 491699 510103 491759
rect 510137 491699 510149 491759
rect 510091 491687 510149 491699
rect 510209 491759 510267 491771
rect 510209 491699 510221 491759
rect 510255 491699 510267 491759
rect 510209 491687 510267 491699
rect 510367 491759 510425 491771
rect 510367 491699 510379 491759
rect 510413 491699 510425 491759
rect 510367 491687 510425 491699
rect 510485 491759 510543 491771
rect 510485 491699 510497 491759
rect 510531 491699 510543 491759
rect 510485 491687 510543 491699
rect 510643 491759 510701 491771
rect 510643 491699 510655 491759
rect 510689 491699 510701 491759
rect 510643 491687 510701 491699
rect 510761 491759 510819 491771
rect 510761 491699 510773 491759
rect 510807 491699 510819 491759
rect 510761 491687 510819 491699
rect 510919 491759 510977 491771
rect 510919 491699 510931 491759
rect 510965 491699 510977 491759
rect 510919 491687 510977 491699
rect 511037 491759 511095 491771
rect 511037 491699 511049 491759
rect 511083 491699 511095 491759
rect 511037 491687 511095 491699
rect 511195 491759 511253 491771
rect 511195 491699 511207 491759
rect 511241 491699 511253 491759
rect 511195 491687 511253 491699
rect 511313 491759 511371 491771
rect 511313 491699 511325 491759
rect 511359 491699 511371 491759
rect 511313 491687 511371 491699
rect 511471 491759 511529 491771
rect 511471 491699 511483 491759
rect 511517 491699 511529 491759
rect 511471 491687 511529 491699
rect 232636 490873 232694 490885
rect 232636 490813 232648 490873
rect 232682 490813 232694 490873
rect 232636 490801 232694 490813
rect 232794 490873 232852 490885
rect 232794 490813 232806 490873
rect 232840 490813 232852 490873
rect 232794 490801 232852 490813
rect 232912 490873 232970 490885
rect 232912 490813 232924 490873
rect 232958 490813 232970 490873
rect 232912 490801 232970 490813
rect 233070 490873 233128 490885
rect 233070 490813 233082 490873
rect 233116 490813 233128 490873
rect 233070 490801 233128 490813
rect 233188 490873 233246 490885
rect 233188 490813 233200 490873
rect 233234 490813 233246 490873
rect 233188 490801 233246 490813
rect 233346 490873 233404 490885
rect 233346 490813 233358 490873
rect 233392 490813 233404 490873
rect 233346 490801 233404 490813
rect 233464 490873 233522 490885
rect 233464 490813 233476 490873
rect 233510 490813 233522 490873
rect 233464 490801 233522 490813
rect 233622 490873 233680 490885
rect 233622 490813 233634 490873
rect 233668 490813 233680 490873
rect 233622 490801 233680 490813
rect 233740 490873 233798 490885
rect 233740 490813 233752 490873
rect 233786 490813 233798 490873
rect 233740 490801 233798 490813
rect 233898 490873 233956 490885
rect 233898 490813 233910 490873
rect 233944 490813 233956 490873
rect 233898 490801 233956 490813
rect 234016 490873 234074 490885
rect 234016 490813 234028 490873
rect 234062 490813 234074 490873
rect 234016 490801 234074 490813
rect 234174 490873 234232 490885
rect 234174 490813 234186 490873
rect 234220 490813 234232 490873
rect 234174 490801 234232 490813
rect 234292 490873 234350 490885
rect 234292 490813 234304 490873
rect 234338 490813 234350 490873
rect 234292 490801 234350 490813
rect 234450 490873 234508 490885
rect 234450 490813 234462 490873
rect 234496 490813 234508 490873
rect 234450 490801 234508 490813
rect 234568 490873 234626 490885
rect 234568 490813 234580 490873
rect 234614 490813 234626 490873
rect 234568 490801 234626 490813
rect 234726 490873 234784 490885
rect 234726 490813 234738 490873
rect 234772 490813 234784 490873
rect 234726 490801 234784 490813
rect 234844 490873 234902 490885
rect 234844 490813 234856 490873
rect 234890 490813 234902 490873
rect 234844 490801 234902 490813
rect 235002 490873 235060 490885
rect 235002 490813 235014 490873
rect 235048 490813 235060 490873
rect 235002 490801 235060 490813
rect 235120 490873 235178 490885
rect 235120 490813 235132 490873
rect 235166 490813 235178 490873
rect 235120 490801 235178 490813
rect 235278 490873 235336 490885
rect 235278 490813 235290 490873
rect 235324 490813 235336 490873
rect 235278 490801 235336 490813
rect 235396 490873 235454 490885
rect 235396 490813 235408 490873
rect 235442 490813 235454 490873
rect 235396 490801 235454 490813
rect 235554 490873 235612 490885
rect 235554 490813 235566 490873
rect 235600 490813 235612 490873
rect 235554 490801 235612 490813
rect 235672 490873 235730 490885
rect 235672 490813 235684 490873
rect 235718 490813 235730 490873
rect 235672 490801 235730 490813
rect 235830 490873 235888 490885
rect 235830 490813 235842 490873
rect 235876 490813 235888 490873
rect 235830 490801 235888 490813
rect 235948 490873 236006 490885
rect 235948 490813 235960 490873
rect 235994 490813 236006 490873
rect 235948 490801 236006 490813
rect 236106 490873 236164 490885
rect 236106 490813 236118 490873
rect 236152 490813 236164 490873
rect 236106 490801 236164 490813
rect 236224 490873 236282 490885
rect 236224 490813 236236 490873
rect 236270 490813 236282 490873
rect 236224 490801 236282 490813
rect 236382 490873 236440 490885
rect 236382 490813 236394 490873
rect 236428 490813 236440 490873
rect 236382 490801 236440 490813
rect 236500 490873 236558 490885
rect 236500 490813 236512 490873
rect 236546 490813 236558 490873
rect 236500 490801 236558 490813
rect 236658 490873 236716 490885
rect 236658 490813 236670 490873
rect 236704 490813 236716 490873
rect 236658 490801 236716 490813
rect 236776 490873 236834 490885
rect 236776 490813 236788 490873
rect 236822 490813 236834 490873
rect 236776 490801 236834 490813
rect 236934 490873 236992 490885
rect 236934 490813 236946 490873
rect 236980 490813 236992 490873
rect 236934 490801 236992 490813
rect 237052 490873 237110 490885
rect 237052 490813 237064 490873
rect 237098 490813 237110 490873
rect 237052 490801 237110 490813
rect 237210 490873 237268 490885
rect 237210 490813 237222 490873
rect 237256 490813 237268 490873
rect 237210 490801 237268 490813
rect 237328 490873 237386 490885
rect 237328 490813 237340 490873
rect 237374 490813 237386 490873
rect 237328 490801 237386 490813
rect 237486 490873 237544 490885
rect 237486 490813 237498 490873
rect 237532 490813 237544 490873
rect 237486 490801 237544 490813
rect 237604 490873 237662 490885
rect 237604 490813 237616 490873
rect 237650 490813 237662 490873
rect 237604 490801 237662 490813
rect 237762 490873 237820 490885
rect 237762 490813 237774 490873
rect 237808 490813 237820 490873
rect 237762 490801 237820 490813
rect 237880 490873 237938 490885
rect 237880 490813 237892 490873
rect 237926 490813 237938 490873
rect 237880 490801 237938 490813
rect 238038 490873 238096 490885
rect 238038 490813 238050 490873
rect 238084 490813 238096 490873
rect 238038 490801 238096 490813
rect 238156 490873 238214 490885
rect 238156 490813 238168 490873
rect 238202 490813 238214 490873
rect 238156 490801 238214 490813
rect 238314 490873 238372 490885
rect 238314 490813 238326 490873
rect 238360 490813 238372 490873
rect 238314 490801 238372 490813
rect 238432 490873 238490 490885
rect 238432 490813 238444 490873
rect 238478 490813 238490 490873
rect 238432 490801 238490 490813
rect 238590 490873 238648 490885
rect 238590 490813 238602 490873
rect 238636 490813 238648 490873
rect 238590 490801 238648 490813
rect 238708 490873 238766 490885
rect 238708 490813 238720 490873
rect 238754 490813 238766 490873
rect 238708 490801 238766 490813
rect 238866 490873 238924 490885
rect 238866 490813 238878 490873
rect 238912 490813 238924 490873
rect 238866 490801 238924 490813
rect 238984 490873 239042 490885
rect 238984 490813 238996 490873
rect 239030 490813 239042 490873
rect 238984 490801 239042 490813
rect 239142 490873 239200 490885
rect 239142 490813 239154 490873
rect 239188 490813 239200 490873
rect 239142 490801 239200 490813
rect 239260 490873 239318 490885
rect 239260 490813 239272 490873
rect 239306 490813 239318 490873
rect 239260 490801 239318 490813
rect 239418 490873 239476 490885
rect 239418 490813 239430 490873
rect 239464 490813 239476 490873
rect 239418 490801 239476 490813
rect 239536 490873 239594 490885
rect 239536 490813 239548 490873
rect 239582 490813 239594 490873
rect 239536 490801 239594 490813
rect 239694 490873 239752 490885
rect 239694 490813 239706 490873
rect 239740 490813 239752 490873
rect 239694 490801 239752 490813
rect 239812 490873 239870 490885
rect 239812 490813 239824 490873
rect 239858 490813 239870 490873
rect 239812 490801 239870 490813
rect 239970 490873 240028 490885
rect 239970 490813 239982 490873
rect 240016 490813 240028 490873
rect 239970 490801 240028 490813
rect 240088 490873 240146 490885
rect 240088 490813 240100 490873
rect 240134 490813 240146 490873
rect 240088 490801 240146 490813
rect 240246 490873 240304 490885
rect 240246 490813 240258 490873
rect 240292 490813 240304 490873
rect 240246 490801 240304 490813
rect 240364 490873 240422 490885
rect 240364 490813 240376 490873
rect 240410 490813 240422 490873
rect 240364 490801 240422 490813
rect 240522 490873 240580 490885
rect 240522 490813 240534 490873
rect 240568 490813 240580 490873
rect 240522 490801 240580 490813
rect 240640 490873 240698 490885
rect 240640 490813 240652 490873
rect 240686 490813 240698 490873
rect 240640 490801 240698 490813
rect 240798 490873 240856 490885
rect 240798 490813 240810 490873
rect 240844 490813 240856 490873
rect 240798 490801 240856 490813
rect 240916 490873 240974 490885
rect 240916 490813 240928 490873
rect 240962 490813 240974 490873
rect 240916 490801 240974 490813
rect 241074 490873 241132 490885
rect 241074 490813 241086 490873
rect 241120 490813 241132 490873
rect 241074 490801 241132 490813
rect 241192 490873 241250 490885
rect 241192 490813 241204 490873
rect 241238 490813 241250 490873
rect 241192 490801 241250 490813
rect 241350 490873 241408 490885
rect 241350 490813 241362 490873
rect 241396 490813 241408 490873
rect 241350 490801 241408 490813
rect 241468 490873 241526 490885
rect 241468 490813 241480 490873
rect 241514 490813 241526 490873
rect 241468 490801 241526 490813
rect 241626 490873 241684 490885
rect 241626 490813 241638 490873
rect 241672 490813 241684 490873
rect 241626 490801 241684 490813
rect 241744 490873 241802 490885
rect 241744 490813 241756 490873
rect 241790 490813 241802 490873
rect 241744 490801 241802 490813
rect 241902 490873 241960 490885
rect 241902 490813 241914 490873
rect 241948 490813 241960 490873
rect 241902 490801 241960 490813
rect 242020 490873 242078 490885
rect 242020 490813 242032 490873
rect 242066 490813 242078 490873
rect 242020 490801 242078 490813
rect 242178 490873 242236 490885
rect 242178 490813 242190 490873
rect 242224 490813 242236 490873
rect 242178 490801 242236 490813
rect 242296 490873 242354 490885
rect 242296 490813 242308 490873
rect 242342 490813 242354 490873
rect 242296 490801 242354 490813
rect 242454 490873 242512 490885
rect 242454 490813 242466 490873
rect 242500 490813 242512 490873
rect 242454 490801 242512 490813
rect 242572 490873 242630 490885
rect 242572 490813 242584 490873
rect 242618 490813 242630 490873
rect 242572 490801 242630 490813
rect 242730 490873 242788 490885
rect 242730 490813 242742 490873
rect 242776 490813 242788 490873
rect 242730 490801 242788 490813
rect 242848 490873 242906 490885
rect 242848 490813 242860 490873
rect 242894 490813 242906 490873
rect 242848 490801 242906 490813
rect 243006 490873 243064 490885
rect 243006 490813 243018 490873
rect 243052 490813 243064 490873
rect 243006 490801 243064 490813
rect 243124 490873 243182 490885
rect 243124 490813 243136 490873
rect 243170 490813 243182 490873
rect 243124 490801 243182 490813
rect 243282 490873 243340 490885
rect 243282 490813 243294 490873
rect 243328 490813 243340 490873
rect 243282 490801 243340 490813
rect 243400 490873 243458 490885
rect 243400 490813 243412 490873
rect 243446 490813 243458 490873
rect 243400 490801 243458 490813
rect 243558 490873 243616 490885
rect 243558 490813 243570 490873
rect 243604 490813 243616 490873
rect 243558 490801 243616 490813
rect 243676 490873 243734 490885
rect 243676 490813 243688 490873
rect 243722 490813 243734 490873
rect 243676 490801 243734 490813
rect 243834 490873 243892 490885
rect 243834 490813 243846 490873
rect 243880 490813 243892 490873
rect 243834 490801 243892 490813
rect 243952 490873 244010 490885
rect 243952 490813 243964 490873
rect 243998 490813 244010 490873
rect 243952 490801 244010 490813
rect 244110 490873 244168 490885
rect 244110 490813 244122 490873
rect 244156 490813 244168 490873
rect 244110 490801 244168 490813
rect 244228 490873 244286 490885
rect 244228 490813 244240 490873
rect 244274 490813 244286 490873
rect 244228 490801 244286 490813
rect 244386 490873 244444 490885
rect 244386 490813 244398 490873
rect 244432 490813 244444 490873
rect 244386 490801 244444 490813
rect 244504 490873 244562 490885
rect 244504 490813 244516 490873
rect 244550 490813 244562 490873
rect 244504 490801 244562 490813
rect 244662 490873 244720 490885
rect 244662 490813 244674 490873
rect 244708 490813 244720 490873
rect 244662 490801 244720 490813
rect 244780 490873 244838 490885
rect 244780 490813 244792 490873
rect 244826 490813 244838 490873
rect 244780 490801 244838 490813
rect 244938 490873 244996 490885
rect 244938 490813 244950 490873
rect 244984 490813 244996 490873
rect 244938 490801 244996 490813
rect 245056 490873 245114 490885
rect 245056 490813 245068 490873
rect 245102 490813 245114 490873
rect 245056 490801 245114 490813
rect 245214 490873 245272 490885
rect 245214 490813 245226 490873
rect 245260 490813 245272 490873
rect 245214 490801 245272 490813
rect 245332 490873 245390 490885
rect 245332 490813 245344 490873
rect 245378 490813 245390 490873
rect 245332 490801 245390 490813
rect 245490 490873 245548 490885
rect 245490 490813 245502 490873
rect 245536 490813 245548 490873
rect 245490 490801 245548 490813
rect 245608 490873 245666 490885
rect 245608 490813 245620 490873
rect 245654 490813 245666 490873
rect 245608 490801 245666 490813
rect 245766 490873 245824 490885
rect 245766 490813 245778 490873
rect 245812 490813 245824 490873
rect 245766 490801 245824 490813
rect 245884 490873 245942 490885
rect 245884 490813 245896 490873
rect 245930 490813 245942 490873
rect 245884 490801 245942 490813
rect 246042 490873 246100 490885
rect 246042 490813 246054 490873
rect 246088 490813 246100 490873
rect 246042 490801 246100 490813
rect 246160 490873 246218 490885
rect 246160 490813 246172 490873
rect 246206 490813 246218 490873
rect 246160 490801 246218 490813
rect 246318 490873 246376 490885
rect 246318 490813 246330 490873
rect 246364 490813 246376 490873
rect 246318 490801 246376 490813
rect 246436 490873 246494 490885
rect 246436 490813 246448 490873
rect 246482 490813 246494 490873
rect 246436 490801 246494 490813
rect 246594 490873 246652 490885
rect 246594 490813 246606 490873
rect 246640 490813 246652 490873
rect 246594 490801 246652 490813
rect 323819 372147 323877 372159
rect 323819 372087 323831 372147
rect 323865 372087 323877 372147
rect 323819 372075 323877 372087
rect 323977 372147 324035 372159
rect 323977 372087 323989 372147
rect 324023 372087 324035 372147
rect 323977 372075 324035 372087
rect 324095 372147 324153 372159
rect 324095 372087 324107 372147
rect 324141 372087 324153 372147
rect 324095 372075 324153 372087
rect 324253 372147 324311 372159
rect 324253 372087 324265 372147
rect 324299 372087 324311 372147
rect 324253 372075 324311 372087
rect 324371 372147 324429 372159
rect 324371 372087 324383 372147
rect 324417 372087 324429 372147
rect 324371 372075 324429 372087
rect 324529 372147 324587 372159
rect 324529 372087 324541 372147
rect 324575 372087 324587 372147
rect 324529 372075 324587 372087
rect 324647 372147 324705 372159
rect 324647 372087 324659 372147
rect 324693 372087 324705 372147
rect 324647 372075 324705 372087
rect 324805 372147 324863 372159
rect 324805 372087 324817 372147
rect 324851 372087 324863 372147
rect 324805 372075 324863 372087
rect 324923 372147 324981 372159
rect 324923 372087 324935 372147
rect 324969 372087 324981 372147
rect 324923 372075 324981 372087
rect 325081 372147 325139 372159
rect 325081 372087 325093 372147
rect 325127 372087 325139 372147
rect 325081 372075 325139 372087
rect 325199 372147 325257 372159
rect 325199 372087 325211 372147
rect 325245 372087 325257 372147
rect 325199 372075 325257 372087
rect 325357 372147 325415 372159
rect 325357 372087 325369 372147
rect 325403 372087 325415 372147
rect 325357 372075 325415 372087
rect 325475 372147 325533 372159
rect 325475 372087 325487 372147
rect 325521 372087 325533 372147
rect 325475 372075 325533 372087
rect 325633 372147 325691 372159
rect 325633 372087 325645 372147
rect 325679 372087 325691 372147
rect 325633 372075 325691 372087
rect 325751 372147 325809 372159
rect 325751 372087 325763 372147
rect 325797 372087 325809 372147
rect 325751 372075 325809 372087
rect 325909 372147 325967 372159
rect 325909 372087 325921 372147
rect 325955 372087 325967 372147
rect 325909 372075 325967 372087
rect 326027 372147 326085 372159
rect 326027 372087 326039 372147
rect 326073 372087 326085 372147
rect 326027 372075 326085 372087
rect 326185 372147 326243 372159
rect 326185 372087 326197 372147
rect 326231 372087 326243 372147
rect 326185 372075 326243 372087
rect 326303 372147 326361 372159
rect 326303 372087 326315 372147
rect 326349 372087 326361 372147
rect 326303 372075 326361 372087
rect 326461 372147 326519 372159
rect 326461 372087 326473 372147
rect 326507 372087 326519 372147
rect 326461 372075 326519 372087
rect 326579 372147 326637 372159
rect 326579 372087 326591 372147
rect 326625 372087 326637 372147
rect 326579 372075 326637 372087
rect 326737 372147 326795 372159
rect 326737 372087 326749 372147
rect 326783 372087 326795 372147
rect 326737 372075 326795 372087
rect 326855 372147 326913 372159
rect 326855 372087 326867 372147
rect 326901 372087 326913 372147
rect 326855 372075 326913 372087
rect 327013 372147 327071 372159
rect 327013 372087 327025 372147
rect 327059 372087 327071 372147
rect 327013 372075 327071 372087
rect 327131 372147 327189 372159
rect 327131 372087 327143 372147
rect 327177 372087 327189 372147
rect 327131 372075 327189 372087
rect 327289 372147 327347 372159
rect 327289 372087 327301 372147
rect 327335 372087 327347 372147
rect 327289 372075 327347 372087
rect 327407 372147 327465 372159
rect 327407 372087 327419 372147
rect 327453 372087 327465 372147
rect 327407 372075 327465 372087
rect 327565 372147 327623 372159
rect 327565 372087 327577 372147
rect 327611 372087 327623 372147
rect 327565 372075 327623 372087
rect 327683 372147 327741 372159
rect 327683 372087 327695 372147
rect 327729 372087 327741 372147
rect 327683 372075 327741 372087
rect 327841 372147 327899 372159
rect 327841 372087 327853 372147
rect 327887 372087 327899 372147
rect 327841 372075 327899 372087
rect 327959 372147 328017 372159
rect 327959 372087 327971 372147
rect 328005 372087 328017 372147
rect 327959 372075 328017 372087
rect 328117 372147 328175 372159
rect 328117 372087 328129 372147
rect 328163 372087 328175 372147
rect 328117 372075 328175 372087
rect 328235 372147 328293 372159
rect 328235 372087 328247 372147
rect 328281 372087 328293 372147
rect 328235 372075 328293 372087
rect 328393 372147 328451 372159
rect 328393 372087 328405 372147
rect 328439 372087 328451 372147
rect 328393 372075 328451 372087
rect 328511 372147 328569 372159
rect 328511 372087 328523 372147
rect 328557 372087 328569 372147
rect 328511 372075 328569 372087
rect 328669 372147 328727 372159
rect 328669 372087 328681 372147
rect 328715 372087 328727 372147
rect 328669 372075 328727 372087
rect 328787 372147 328845 372159
rect 328787 372087 328799 372147
rect 328833 372087 328845 372147
rect 328787 372075 328845 372087
rect 328945 372147 329003 372159
rect 328945 372087 328957 372147
rect 328991 372087 329003 372147
rect 328945 372075 329003 372087
rect 329063 372147 329121 372159
rect 329063 372087 329075 372147
rect 329109 372087 329121 372147
rect 329063 372075 329121 372087
rect 329221 372147 329279 372159
rect 329221 372087 329233 372147
rect 329267 372087 329279 372147
rect 329221 372075 329279 372087
rect 329339 372147 329397 372159
rect 329339 372087 329351 372147
rect 329385 372087 329397 372147
rect 329339 372075 329397 372087
rect 329497 372147 329555 372159
rect 329497 372087 329509 372147
rect 329543 372087 329555 372147
rect 329497 372075 329555 372087
rect 329615 372147 329673 372159
rect 329615 372087 329627 372147
rect 329661 372087 329673 372147
rect 329615 372075 329673 372087
rect 329773 372147 329831 372159
rect 329773 372087 329785 372147
rect 329819 372087 329831 372147
rect 329773 372075 329831 372087
rect 329891 372147 329949 372159
rect 329891 372087 329903 372147
rect 329937 372087 329949 372147
rect 329891 372075 329949 372087
rect 330049 372147 330107 372159
rect 330049 372087 330061 372147
rect 330095 372087 330107 372147
rect 330049 372075 330107 372087
rect 330167 372147 330225 372159
rect 330167 372087 330179 372147
rect 330213 372087 330225 372147
rect 330167 372075 330225 372087
rect 330325 372147 330383 372159
rect 330325 372087 330337 372147
rect 330371 372087 330383 372147
rect 330325 372075 330383 372087
rect 330443 372147 330501 372159
rect 330443 372087 330455 372147
rect 330489 372087 330501 372147
rect 330443 372075 330501 372087
rect 330601 372147 330659 372159
rect 330601 372087 330613 372147
rect 330647 372087 330659 372147
rect 330601 372075 330659 372087
rect 330719 372147 330777 372159
rect 330719 372087 330731 372147
rect 330765 372087 330777 372147
rect 330719 372075 330777 372087
rect 330877 372147 330935 372159
rect 330877 372087 330889 372147
rect 330923 372087 330935 372147
rect 330877 372075 330935 372087
rect 330995 372147 331053 372159
rect 330995 372087 331007 372147
rect 331041 372087 331053 372147
rect 330995 372075 331053 372087
rect 331153 372147 331211 372159
rect 331153 372087 331165 372147
rect 331199 372087 331211 372147
rect 331153 372075 331211 372087
rect 331271 372147 331329 372159
rect 331271 372087 331283 372147
rect 331317 372087 331329 372147
rect 331271 372075 331329 372087
rect 331429 372147 331487 372159
rect 331429 372087 331441 372147
rect 331475 372087 331487 372147
rect 331429 372075 331487 372087
rect 331547 372147 331605 372159
rect 331547 372087 331559 372147
rect 331593 372087 331605 372147
rect 331547 372075 331605 372087
rect 331705 372147 331763 372159
rect 331705 372087 331717 372147
rect 331751 372087 331763 372147
rect 331705 372075 331763 372087
rect 331823 372147 331881 372159
rect 331823 372087 331835 372147
rect 331869 372087 331881 372147
rect 331823 372075 331881 372087
rect 331981 372147 332039 372159
rect 331981 372087 331993 372147
rect 332027 372087 332039 372147
rect 331981 372075 332039 372087
rect 332099 372147 332157 372159
rect 332099 372087 332111 372147
rect 332145 372087 332157 372147
rect 332099 372075 332157 372087
rect 332257 372147 332315 372159
rect 332257 372087 332269 372147
rect 332303 372087 332315 372147
rect 332257 372075 332315 372087
rect 332375 372147 332433 372159
rect 332375 372087 332387 372147
rect 332421 372087 332433 372147
rect 332375 372075 332433 372087
rect 332533 372147 332591 372159
rect 332533 372087 332545 372147
rect 332579 372087 332591 372147
rect 332533 372075 332591 372087
rect 332651 372147 332709 372159
rect 332651 372087 332663 372147
rect 332697 372087 332709 372147
rect 332651 372075 332709 372087
rect 332809 372147 332867 372159
rect 332809 372087 332821 372147
rect 332855 372087 332867 372147
rect 332809 372075 332867 372087
rect 332927 372147 332985 372159
rect 332927 372087 332939 372147
rect 332973 372087 332985 372147
rect 332927 372075 332985 372087
rect 333085 372147 333143 372159
rect 333085 372087 333097 372147
rect 333131 372087 333143 372147
rect 333085 372075 333143 372087
rect 333203 372147 333261 372159
rect 333203 372087 333215 372147
rect 333249 372087 333261 372147
rect 333203 372075 333261 372087
rect 333361 372147 333419 372159
rect 333361 372087 333373 372147
rect 333407 372087 333419 372147
rect 333361 372075 333419 372087
rect 333479 372147 333537 372159
rect 333479 372087 333491 372147
rect 333525 372087 333537 372147
rect 333479 372075 333537 372087
rect 333637 372147 333695 372159
rect 333637 372087 333649 372147
rect 333683 372087 333695 372147
rect 333637 372075 333695 372087
rect 333755 372147 333813 372159
rect 333755 372087 333767 372147
rect 333801 372087 333813 372147
rect 333755 372075 333813 372087
rect 333913 372147 333971 372159
rect 333913 372087 333925 372147
rect 333959 372087 333971 372147
rect 333913 372075 333971 372087
rect 334031 372147 334089 372159
rect 334031 372087 334043 372147
rect 334077 372087 334089 372147
rect 334031 372075 334089 372087
rect 334189 372147 334247 372159
rect 334189 372087 334201 372147
rect 334235 372087 334247 372147
rect 334189 372075 334247 372087
rect 334307 372147 334365 372159
rect 334307 372087 334319 372147
rect 334353 372087 334365 372147
rect 334307 372075 334365 372087
rect 334465 372147 334523 372159
rect 334465 372087 334477 372147
rect 334511 372087 334523 372147
rect 334465 372075 334523 372087
rect 334583 372147 334641 372159
rect 334583 372087 334595 372147
rect 334629 372087 334641 372147
rect 334583 372075 334641 372087
rect 334741 372147 334799 372159
rect 334741 372087 334753 372147
rect 334787 372087 334799 372147
rect 334741 372075 334799 372087
rect 334859 372147 334917 372159
rect 334859 372087 334871 372147
rect 334905 372087 334917 372147
rect 334859 372075 334917 372087
rect 335017 372147 335075 372159
rect 335017 372087 335029 372147
rect 335063 372087 335075 372147
rect 335017 372075 335075 372087
rect 335135 372147 335193 372159
rect 335135 372087 335147 372147
rect 335181 372087 335193 372147
rect 335135 372075 335193 372087
rect 335293 372147 335351 372159
rect 335293 372087 335305 372147
rect 335339 372087 335351 372147
rect 335293 372075 335351 372087
rect 335411 372147 335469 372159
rect 335411 372087 335423 372147
rect 335457 372087 335469 372147
rect 335411 372075 335469 372087
rect 335569 372147 335627 372159
rect 335569 372087 335581 372147
rect 335615 372087 335627 372147
rect 335569 372075 335627 372087
rect 335687 372147 335745 372159
rect 335687 372087 335699 372147
rect 335733 372087 335745 372147
rect 335687 372075 335745 372087
rect 335845 372147 335903 372159
rect 335845 372087 335857 372147
rect 335891 372087 335903 372147
rect 335845 372075 335903 372087
rect 335963 372147 336021 372159
rect 335963 372087 335975 372147
rect 336009 372087 336021 372147
rect 335963 372075 336021 372087
rect 336121 372147 336179 372159
rect 336121 372087 336133 372147
rect 336167 372087 336179 372147
rect 336121 372075 336179 372087
rect 336239 372147 336297 372159
rect 336239 372087 336251 372147
rect 336285 372087 336297 372147
rect 336239 372075 336297 372087
rect 336397 372147 336455 372159
rect 336397 372087 336409 372147
rect 336443 372087 336455 372147
rect 336397 372075 336455 372087
rect 336515 372147 336573 372159
rect 336515 372087 336527 372147
rect 336561 372087 336573 372147
rect 336515 372075 336573 372087
rect 336673 372147 336731 372159
rect 336673 372087 336685 372147
rect 336719 372087 336731 372147
rect 336673 372075 336731 372087
rect 336791 372147 336849 372159
rect 336791 372087 336803 372147
rect 336837 372087 336849 372147
rect 336791 372075 336849 372087
rect 336949 372147 337007 372159
rect 336949 372087 336961 372147
rect 336995 372087 337007 372147
rect 336949 372075 337007 372087
rect 337067 372147 337125 372159
rect 337067 372087 337079 372147
rect 337113 372087 337125 372147
rect 337067 372075 337125 372087
rect 337225 372147 337283 372159
rect 337225 372087 337237 372147
rect 337271 372087 337283 372147
rect 337225 372075 337283 372087
rect 337343 372147 337401 372159
rect 337343 372087 337355 372147
rect 337389 372087 337401 372147
rect 337343 372075 337401 372087
rect 337501 372147 337559 372159
rect 337501 372087 337513 372147
rect 337547 372087 337559 372147
rect 337501 372075 337559 372087
rect 337619 372147 337677 372159
rect 337619 372087 337631 372147
rect 337665 372087 337677 372147
rect 337619 372075 337677 372087
rect 337777 372147 337835 372159
rect 337777 372087 337789 372147
rect 337823 372087 337835 372147
rect 337777 372075 337835 372087
rect 53279 371469 53337 371481
rect 53279 371409 53291 371469
rect 53325 371409 53337 371469
rect 53279 371397 53337 371409
rect 53437 371469 53495 371481
rect 53437 371409 53449 371469
rect 53483 371409 53495 371469
rect 53437 371397 53495 371409
rect 53555 371469 53613 371481
rect 53555 371409 53567 371469
rect 53601 371409 53613 371469
rect 53555 371397 53613 371409
rect 53713 371469 53771 371481
rect 53713 371409 53725 371469
rect 53759 371409 53771 371469
rect 53713 371397 53771 371409
rect 53831 371469 53889 371481
rect 53831 371409 53843 371469
rect 53877 371409 53889 371469
rect 53831 371397 53889 371409
rect 53989 371469 54047 371481
rect 53989 371409 54001 371469
rect 54035 371409 54047 371469
rect 53989 371397 54047 371409
rect 54107 371469 54165 371481
rect 54107 371409 54119 371469
rect 54153 371409 54165 371469
rect 54107 371397 54165 371409
rect 54265 371469 54323 371481
rect 54265 371409 54277 371469
rect 54311 371409 54323 371469
rect 54265 371397 54323 371409
rect 54383 371469 54441 371481
rect 54383 371409 54395 371469
rect 54429 371409 54441 371469
rect 54383 371397 54441 371409
rect 54541 371469 54599 371481
rect 54541 371409 54553 371469
rect 54587 371409 54599 371469
rect 54541 371397 54599 371409
rect 54659 371469 54717 371481
rect 54659 371409 54671 371469
rect 54705 371409 54717 371469
rect 54659 371397 54717 371409
rect 54817 371469 54875 371481
rect 54817 371409 54829 371469
rect 54863 371409 54875 371469
rect 54817 371397 54875 371409
rect 54935 371469 54993 371481
rect 54935 371409 54947 371469
rect 54981 371409 54993 371469
rect 54935 371397 54993 371409
rect 55093 371469 55151 371481
rect 55093 371409 55105 371469
rect 55139 371409 55151 371469
rect 55093 371397 55151 371409
rect 55211 371469 55269 371481
rect 55211 371409 55223 371469
rect 55257 371409 55269 371469
rect 55211 371397 55269 371409
rect 55369 371469 55427 371481
rect 55369 371409 55381 371469
rect 55415 371409 55427 371469
rect 55369 371397 55427 371409
rect 55487 371469 55545 371481
rect 55487 371409 55499 371469
rect 55533 371409 55545 371469
rect 55487 371397 55545 371409
rect 55645 371469 55703 371481
rect 55645 371409 55657 371469
rect 55691 371409 55703 371469
rect 55645 371397 55703 371409
rect 55763 371469 55821 371481
rect 55763 371409 55775 371469
rect 55809 371409 55821 371469
rect 55763 371397 55821 371409
rect 55921 371469 55979 371481
rect 55921 371409 55933 371469
rect 55967 371409 55979 371469
rect 55921 371397 55979 371409
rect 56039 371469 56097 371481
rect 56039 371409 56051 371469
rect 56085 371409 56097 371469
rect 56039 371397 56097 371409
rect 56197 371469 56255 371481
rect 56197 371409 56209 371469
rect 56243 371409 56255 371469
rect 56197 371397 56255 371409
rect 56315 371469 56373 371481
rect 56315 371409 56327 371469
rect 56361 371409 56373 371469
rect 56315 371397 56373 371409
rect 56473 371469 56531 371481
rect 56473 371409 56485 371469
rect 56519 371409 56531 371469
rect 56473 371397 56531 371409
rect 56591 371469 56649 371481
rect 56591 371409 56603 371469
rect 56637 371409 56649 371469
rect 56591 371397 56649 371409
rect 56749 371469 56807 371481
rect 56749 371409 56761 371469
rect 56795 371409 56807 371469
rect 56749 371397 56807 371409
rect 56867 371469 56925 371481
rect 56867 371409 56879 371469
rect 56913 371409 56925 371469
rect 56867 371397 56925 371409
rect 57025 371469 57083 371481
rect 57025 371409 57037 371469
rect 57071 371409 57083 371469
rect 57025 371397 57083 371409
rect 57143 371469 57201 371481
rect 57143 371409 57155 371469
rect 57189 371409 57201 371469
rect 57143 371397 57201 371409
rect 57301 371469 57359 371481
rect 57301 371409 57313 371469
rect 57347 371409 57359 371469
rect 57301 371397 57359 371409
rect 57419 371469 57477 371481
rect 57419 371409 57431 371469
rect 57465 371409 57477 371469
rect 57419 371397 57477 371409
rect 57577 371469 57635 371481
rect 57577 371409 57589 371469
rect 57623 371409 57635 371469
rect 57577 371397 57635 371409
rect 57695 371469 57753 371481
rect 57695 371409 57707 371469
rect 57741 371409 57753 371469
rect 57695 371397 57753 371409
rect 57853 371469 57911 371481
rect 57853 371409 57865 371469
rect 57899 371409 57911 371469
rect 57853 371397 57911 371409
rect 57971 371469 58029 371481
rect 57971 371409 57983 371469
rect 58017 371409 58029 371469
rect 57971 371397 58029 371409
rect 58129 371469 58187 371481
rect 58129 371409 58141 371469
rect 58175 371409 58187 371469
rect 58129 371397 58187 371409
rect 58247 371469 58305 371481
rect 58247 371409 58259 371469
rect 58293 371409 58305 371469
rect 58247 371397 58305 371409
rect 58405 371469 58463 371481
rect 58405 371409 58417 371469
rect 58451 371409 58463 371469
rect 58405 371397 58463 371409
rect 58523 371469 58581 371481
rect 58523 371409 58535 371469
rect 58569 371409 58581 371469
rect 58523 371397 58581 371409
rect 58681 371469 58739 371481
rect 58681 371409 58693 371469
rect 58727 371409 58739 371469
rect 58681 371397 58739 371409
rect 58799 371469 58857 371481
rect 58799 371409 58811 371469
rect 58845 371409 58857 371469
rect 58799 371397 58857 371409
rect 58957 371469 59015 371481
rect 58957 371409 58969 371469
rect 59003 371409 59015 371469
rect 58957 371397 59015 371409
rect 59075 371469 59133 371481
rect 59075 371409 59087 371469
rect 59121 371409 59133 371469
rect 59075 371397 59133 371409
rect 59233 371469 59291 371481
rect 59233 371409 59245 371469
rect 59279 371409 59291 371469
rect 59233 371397 59291 371409
rect 59351 371469 59409 371481
rect 59351 371409 59363 371469
rect 59397 371409 59409 371469
rect 59351 371397 59409 371409
rect 59509 371469 59567 371481
rect 59509 371409 59521 371469
rect 59555 371409 59567 371469
rect 59509 371397 59567 371409
rect 59627 371469 59685 371481
rect 59627 371409 59639 371469
rect 59673 371409 59685 371469
rect 59627 371397 59685 371409
rect 59785 371469 59843 371481
rect 59785 371409 59797 371469
rect 59831 371409 59843 371469
rect 59785 371397 59843 371409
rect 59903 371469 59961 371481
rect 59903 371409 59915 371469
rect 59949 371409 59961 371469
rect 59903 371397 59961 371409
rect 60061 371469 60119 371481
rect 60061 371409 60073 371469
rect 60107 371409 60119 371469
rect 60061 371397 60119 371409
rect 60179 371469 60237 371481
rect 60179 371409 60191 371469
rect 60225 371409 60237 371469
rect 60179 371397 60237 371409
rect 60337 371469 60395 371481
rect 60337 371409 60349 371469
rect 60383 371409 60395 371469
rect 60337 371397 60395 371409
rect 60455 371469 60513 371481
rect 60455 371409 60467 371469
rect 60501 371409 60513 371469
rect 60455 371397 60513 371409
rect 60613 371469 60671 371481
rect 60613 371409 60625 371469
rect 60659 371409 60671 371469
rect 60613 371397 60671 371409
rect 60731 371469 60789 371481
rect 60731 371409 60743 371469
rect 60777 371409 60789 371469
rect 60731 371397 60789 371409
rect 60889 371469 60947 371481
rect 60889 371409 60901 371469
rect 60935 371409 60947 371469
rect 60889 371397 60947 371409
rect 61007 371469 61065 371481
rect 61007 371409 61019 371469
rect 61053 371409 61065 371469
rect 61007 371397 61065 371409
rect 61165 371469 61223 371481
rect 61165 371409 61177 371469
rect 61211 371409 61223 371469
rect 61165 371397 61223 371409
rect 61283 371469 61341 371481
rect 61283 371409 61295 371469
rect 61329 371409 61341 371469
rect 61283 371397 61341 371409
rect 61441 371469 61499 371481
rect 61441 371409 61453 371469
rect 61487 371409 61499 371469
rect 61441 371397 61499 371409
rect 61559 371469 61617 371481
rect 61559 371409 61571 371469
rect 61605 371409 61617 371469
rect 61559 371397 61617 371409
rect 61717 371469 61775 371481
rect 61717 371409 61729 371469
rect 61763 371409 61775 371469
rect 61717 371397 61775 371409
rect 61835 371469 61893 371481
rect 61835 371409 61847 371469
rect 61881 371409 61893 371469
rect 61835 371397 61893 371409
rect 61993 371469 62051 371481
rect 61993 371409 62005 371469
rect 62039 371409 62051 371469
rect 61993 371397 62051 371409
rect 62111 371469 62169 371481
rect 62111 371409 62123 371469
rect 62157 371409 62169 371469
rect 62111 371397 62169 371409
rect 62269 371469 62327 371481
rect 62269 371409 62281 371469
rect 62315 371409 62327 371469
rect 62269 371397 62327 371409
rect 62387 371469 62445 371481
rect 62387 371409 62399 371469
rect 62433 371409 62445 371469
rect 62387 371397 62445 371409
rect 62545 371469 62603 371481
rect 62545 371409 62557 371469
rect 62591 371409 62603 371469
rect 62545 371397 62603 371409
rect 62663 371469 62721 371481
rect 62663 371409 62675 371469
rect 62709 371409 62721 371469
rect 62663 371397 62721 371409
rect 62821 371469 62879 371481
rect 62821 371409 62833 371469
rect 62867 371409 62879 371469
rect 62821 371397 62879 371409
rect 62939 371469 62997 371481
rect 62939 371409 62951 371469
rect 62985 371409 62997 371469
rect 62939 371397 62997 371409
rect 63097 371469 63155 371481
rect 63097 371409 63109 371469
rect 63143 371409 63155 371469
rect 63097 371397 63155 371409
rect 63215 371469 63273 371481
rect 63215 371409 63227 371469
rect 63261 371409 63273 371469
rect 63215 371397 63273 371409
rect 63373 371469 63431 371481
rect 63373 371409 63385 371469
rect 63419 371409 63431 371469
rect 63373 371397 63431 371409
rect 63491 371469 63549 371481
rect 63491 371409 63503 371469
rect 63537 371409 63549 371469
rect 63491 371397 63549 371409
rect 63649 371469 63707 371481
rect 63649 371409 63661 371469
rect 63695 371409 63707 371469
rect 63649 371397 63707 371409
rect 63767 371469 63825 371481
rect 63767 371409 63779 371469
rect 63813 371409 63825 371469
rect 63767 371397 63825 371409
rect 63925 371469 63983 371481
rect 63925 371409 63937 371469
rect 63971 371409 63983 371469
rect 63925 371397 63983 371409
rect 64043 371469 64101 371481
rect 64043 371409 64055 371469
rect 64089 371409 64101 371469
rect 64043 371397 64101 371409
rect 64201 371469 64259 371481
rect 64201 371409 64213 371469
rect 64247 371409 64259 371469
rect 64201 371397 64259 371409
rect 64319 371469 64377 371481
rect 64319 371409 64331 371469
rect 64365 371409 64377 371469
rect 64319 371397 64377 371409
rect 64477 371469 64535 371481
rect 64477 371409 64489 371469
rect 64523 371409 64535 371469
rect 64477 371397 64535 371409
rect 64595 371469 64653 371481
rect 64595 371409 64607 371469
rect 64641 371409 64653 371469
rect 64595 371397 64653 371409
rect 64753 371469 64811 371481
rect 64753 371409 64765 371469
rect 64799 371409 64811 371469
rect 64753 371397 64811 371409
rect 64871 371469 64929 371481
rect 64871 371409 64883 371469
rect 64917 371409 64929 371469
rect 64871 371397 64929 371409
rect 65029 371469 65087 371481
rect 65029 371409 65041 371469
rect 65075 371409 65087 371469
rect 65029 371397 65087 371409
rect 65147 371469 65205 371481
rect 65147 371409 65159 371469
rect 65193 371409 65205 371469
rect 65147 371397 65205 371409
rect 65305 371469 65363 371481
rect 65305 371409 65317 371469
rect 65351 371409 65363 371469
rect 65305 371397 65363 371409
rect 65423 371469 65481 371481
rect 65423 371409 65435 371469
rect 65469 371409 65481 371469
rect 65423 371397 65481 371409
rect 65581 371469 65639 371481
rect 65581 371409 65593 371469
rect 65627 371409 65639 371469
rect 65581 371397 65639 371409
rect 65699 371469 65757 371481
rect 65699 371409 65711 371469
rect 65745 371409 65757 371469
rect 65699 371397 65757 371409
rect 65857 371469 65915 371481
rect 65857 371409 65869 371469
rect 65903 371409 65915 371469
rect 65857 371397 65915 371409
rect 65975 371469 66033 371481
rect 65975 371409 65987 371469
rect 66021 371409 66033 371469
rect 65975 371397 66033 371409
rect 66133 371469 66191 371481
rect 66133 371409 66145 371469
rect 66179 371409 66191 371469
rect 66133 371397 66191 371409
rect 66251 371469 66309 371481
rect 66251 371409 66263 371469
rect 66297 371409 66309 371469
rect 66251 371397 66309 371409
rect 66409 371469 66467 371481
rect 66409 371409 66421 371469
rect 66455 371409 66467 371469
rect 66409 371397 66467 371409
rect 66527 371469 66585 371481
rect 66527 371409 66539 371469
rect 66573 371409 66585 371469
rect 66527 371397 66585 371409
rect 66685 371469 66743 371481
rect 66685 371409 66697 371469
rect 66731 371409 66743 371469
rect 66685 371397 66743 371409
rect 66803 371469 66861 371481
rect 66803 371409 66815 371469
rect 66849 371409 66861 371469
rect 66803 371397 66861 371409
rect 66961 371469 67019 371481
rect 66961 371409 66973 371469
rect 67007 371409 67019 371469
rect 66961 371397 67019 371409
rect 67079 371469 67137 371481
rect 67079 371409 67091 371469
rect 67125 371409 67137 371469
rect 67079 371397 67137 371409
rect 67237 371469 67295 371481
rect 67237 371409 67249 371469
rect 67283 371409 67295 371469
rect 67237 371397 67295 371409
rect 143279 371469 143337 371481
rect 143279 371409 143291 371469
rect 143325 371409 143337 371469
rect 143279 371397 143337 371409
rect 143437 371469 143495 371481
rect 143437 371409 143449 371469
rect 143483 371409 143495 371469
rect 143437 371397 143495 371409
rect 143555 371469 143613 371481
rect 143555 371409 143567 371469
rect 143601 371409 143613 371469
rect 143555 371397 143613 371409
rect 143713 371469 143771 371481
rect 143713 371409 143725 371469
rect 143759 371409 143771 371469
rect 143713 371397 143771 371409
rect 143831 371469 143889 371481
rect 143831 371409 143843 371469
rect 143877 371409 143889 371469
rect 143831 371397 143889 371409
rect 143989 371469 144047 371481
rect 143989 371409 144001 371469
rect 144035 371409 144047 371469
rect 143989 371397 144047 371409
rect 144107 371469 144165 371481
rect 144107 371409 144119 371469
rect 144153 371409 144165 371469
rect 144107 371397 144165 371409
rect 144265 371469 144323 371481
rect 144265 371409 144277 371469
rect 144311 371409 144323 371469
rect 144265 371397 144323 371409
rect 144383 371469 144441 371481
rect 144383 371409 144395 371469
rect 144429 371409 144441 371469
rect 144383 371397 144441 371409
rect 144541 371469 144599 371481
rect 144541 371409 144553 371469
rect 144587 371409 144599 371469
rect 144541 371397 144599 371409
rect 144659 371469 144717 371481
rect 144659 371409 144671 371469
rect 144705 371409 144717 371469
rect 144659 371397 144717 371409
rect 144817 371469 144875 371481
rect 144817 371409 144829 371469
rect 144863 371409 144875 371469
rect 144817 371397 144875 371409
rect 144935 371469 144993 371481
rect 144935 371409 144947 371469
rect 144981 371409 144993 371469
rect 144935 371397 144993 371409
rect 145093 371469 145151 371481
rect 145093 371409 145105 371469
rect 145139 371409 145151 371469
rect 145093 371397 145151 371409
rect 145211 371469 145269 371481
rect 145211 371409 145223 371469
rect 145257 371409 145269 371469
rect 145211 371397 145269 371409
rect 145369 371469 145427 371481
rect 145369 371409 145381 371469
rect 145415 371409 145427 371469
rect 145369 371397 145427 371409
rect 145487 371469 145545 371481
rect 145487 371409 145499 371469
rect 145533 371409 145545 371469
rect 145487 371397 145545 371409
rect 145645 371469 145703 371481
rect 145645 371409 145657 371469
rect 145691 371409 145703 371469
rect 145645 371397 145703 371409
rect 145763 371469 145821 371481
rect 145763 371409 145775 371469
rect 145809 371409 145821 371469
rect 145763 371397 145821 371409
rect 145921 371469 145979 371481
rect 145921 371409 145933 371469
rect 145967 371409 145979 371469
rect 145921 371397 145979 371409
rect 146039 371469 146097 371481
rect 146039 371409 146051 371469
rect 146085 371409 146097 371469
rect 146039 371397 146097 371409
rect 146197 371469 146255 371481
rect 146197 371409 146209 371469
rect 146243 371409 146255 371469
rect 146197 371397 146255 371409
rect 146315 371469 146373 371481
rect 146315 371409 146327 371469
rect 146361 371409 146373 371469
rect 146315 371397 146373 371409
rect 146473 371469 146531 371481
rect 146473 371409 146485 371469
rect 146519 371409 146531 371469
rect 146473 371397 146531 371409
rect 146591 371469 146649 371481
rect 146591 371409 146603 371469
rect 146637 371409 146649 371469
rect 146591 371397 146649 371409
rect 146749 371469 146807 371481
rect 146749 371409 146761 371469
rect 146795 371409 146807 371469
rect 146749 371397 146807 371409
rect 146867 371469 146925 371481
rect 146867 371409 146879 371469
rect 146913 371409 146925 371469
rect 146867 371397 146925 371409
rect 147025 371469 147083 371481
rect 147025 371409 147037 371469
rect 147071 371409 147083 371469
rect 147025 371397 147083 371409
rect 147143 371469 147201 371481
rect 147143 371409 147155 371469
rect 147189 371409 147201 371469
rect 147143 371397 147201 371409
rect 147301 371469 147359 371481
rect 147301 371409 147313 371469
rect 147347 371409 147359 371469
rect 147301 371397 147359 371409
rect 147419 371469 147477 371481
rect 147419 371409 147431 371469
rect 147465 371409 147477 371469
rect 147419 371397 147477 371409
rect 147577 371469 147635 371481
rect 147577 371409 147589 371469
rect 147623 371409 147635 371469
rect 147577 371397 147635 371409
rect 147695 371469 147753 371481
rect 147695 371409 147707 371469
rect 147741 371409 147753 371469
rect 147695 371397 147753 371409
rect 147853 371469 147911 371481
rect 147853 371409 147865 371469
rect 147899 371409 147911 371469
rect 147853 371397 147911 371409
rect 147971 371469 148029 371481
rect 147971 371409 147983 371469
rect 148017 371409 148029 371469
rect 147971 371397 148029 371409
rect 148129 371469 148187 371481
rect 148129 371409 148141 371469
rect 148175 371409 148187 371469
rect 148129 371397 148187 371409
rect 148247 371469 148305 371481
rect 148247 371409 148259 371469
rect 148293 371409 148305 371469
rect 148247 371397 148305 371409
rect 148405 371469 148463 371481
rect 148405 371409 148417 371469
rect 148451 371409 148463 371469
rect 148405 371397 148463 371409
rect 148523 371469 148581 371481
rect 148523 371409 148535 371469
rect 148569 371409 148581 371469
rect 148523 371397 148581 371409
rect 148681 371469 148739 371481
rect 148681 371409 148693 371469
rect 148727 371409 148739 371469
rect 148681 371397 148739 371409
rect 148799 371469 148857 371481
rect 148799 371409 148811 371469
rect 148845 371409 148857 371469
rect 148799 371397 148857 371409
rect 148957 371469 149015 371481
rect 148957 371409 148969 371469
rect 149003 371409 149015 371469
rect 148957 371397 149015 371409
rect 149075 371469 149133 371481
rect 149075 371409 149087 371469
rect 149121 371409 149133 371469
rect 149075 371397 149133 371409
rect 149233 371469 149291 371481
rect 149233 371409 149245 371469
rect 149279 371409 149291 371469
rect 149233 371397 149291 371409
rect 149351 371469 149409 371481
rect 149351 371409 149363 371469
rect 149397 371409 149409 371469
rect 149351 371397 149409 371409
rect 149509 371469 149567 371481
rect 149509 371409 149521 371469
rect 149555 371409 149567 371469
rect 149509 371397 149567 371409
rect 149627 371469 149685 371481
rect 149627 371409 149639 371469
rect 149673 371409 149685 371469
rect 149627 371397 149685 371409
rect 149785 371469 149843 371481
rect 149785 371409 149797 371469
rect 149831 371409 149843 371469
rect 149785 371397 149843 371409
rect 149903 371469 149961 371481
rect 149903 371409 149915 371469
rect 149949 371409 149961 371469
rect 149903 371397 149961 371409
rect 150061 371469 150119 371481
rect 150061 371409 150073 371469
rect 150107 371409 150119 371469
rect 150061 371397 150119 371409
rect 150179 371469 150237 371481
rect 150179 371409 150191 371469
rect 150225 371409 150237 371469
rect 150179 371397 150237 371409
rect 150337 371469 150395 371481
rect 150337 371409 150349 371469
rect 150383 371409 150395 371469
rect 150337 371397 150395 371409
rect 150455 371469 150513 371481
rect 150455 371409 150467 371469
rect 150501 371409 150513 371469
rect 150455 371397 150513 371409
rect 150613 371469 150671 371481
rect 150613 371409 150625 371469
rect 150659 371409 150671 371469
rect 150613 371397 150671 371409
rect 150731 371469 150789 371481
rect 150731 371409 150743 371469
rect 150777 371409 150789 371469
rect 150731 371397 150789 371409
rect 150889 371469 150947 371481
rect 150889 371409 150901 371469
rect 150935 371409 150947 371469
rect 150889 371397 150947 371409
rect 151007 371469 151065 371481
rect 151007 371409 151019 371469
rect 151053 371409 151065 371469
rect 151007 371397 151065 371409
rect 151165 371469 151223 371481
rect 151165 371409 151177 371469
rect 151211 371409 151223 371469
rect 151165 371397 151223 371409
rect 151283 371469 151341 371481
rect 151283 371409 151295 371469
rect 151329 371409 151341 371469
rect 151283 371397 151341 371409
rect 151441 371469 151499 371481
rect 151441 371409 151453 371469
rect 151487 371409 151499 371469
rect 151441 371397 151499 371409
rect 151559 371469 151617 371481
rect 151559 371409 151571 371469
rect 151605 371409 151617 371469
rect 151559 371397 151617 371409
rect 151717 371469 151775 371481
rect 151717 371409 151729 371469
rect 151763 371409 151775 371469
rect 151717 371397 151775 371409
rect 151835 371469 151893 371481
rect 151835 371409 151847 371469
rect 151881 371409 151893 371469
rect 151835 371397 151893 371409
rect 151993 371469 152051 371481
rect 151993 371409 152005 371469
rect 152039 371409 152051 371469
rect 151993 371397 152051 371409
rect 152111 371469 152169 371481
rect 152111 371409 152123 371469
rect 152157 371409 152169 371469
rect 152111 371397 152169 371409
rect 152269 371469 152327 371481
rect 152269 371409 152281 371469
rect 152315 371409 152327 371469
rect 152269 371397 152327 371409
rect 152387 371469 152445 371481
rect 152387 371409 152399 371469
rect 152433 371409 152445 371469
rect 152387 371397 152445 371409
rect 152545 371469 152603 371481
rect 152545 371409 152557 371469
rect 152591 371409 152603 371469
rect 152545 371397 152603 371409
rect 152663 371469 152721 371481
rect 152663 371409 152675 371469
rect 152709 371409 152721 371469
rect 152663 371397 152721 371409
rect 152821 371469 152879 371481
rect 152821 371409 152833 371469
rect 152867 371409 152879 371469
rect 152821 371397 152879 371409
rect 152939 371469 152997 371481
rect 152939 371409 152951 371469
rect 152985 371409 152997 371469
rect 152939 371397 152997 371409
rect 153097 371469 153155 371481
rect 153097 371409 153109 371469
rect 153143 371409 153155 371469
rect 153097 371397 153155 371409
rect 153215 371469 153273 371481
rect 153215 371409 153227 371469
rect 153261 371409 153273 371469
rect 153215 371397 153273 371409
rect 153373 371469 153431 371481
rect 153373 371409 153385 371469
rect 153419 371409 153431 371469
rect 153373 371397 153431 371409
rect 153491 371469 153549 371481
rect 153491 371409 153503 371469
rect 153537 371409 153549 371469
rect 153491 371397 153549 371409
rect 153649 371469 153707 371481
rect 153649 371409 153661 371469
rect 153695 371409 153707 371469
rect 153649 371397 153707 371409
rect 153767 371469 153825 371481
rect 153767 371409 153779 371469
rect 153813 371409 153825 371469
rect 153767 371397 153825 371409
rect 153925 371469 153983 371481
rect 153925 371409 153937 371469
rect 153971 371409 153983 371469
rect 153925 371397 153983 371409
rect 154043 371469 154101 371481
rect 154043 371409 154055 371469
rect 154089 371409 154101 371469
rect 154043 371397 154101 371409
rect 154201 371469 154259 371481
rect 154201 371409 154213 371469
rect 154247 371409 154259 371469
rect 154201 371397 154259 371409
rect 154319 371469 154377 371481
rect 154319 371409 154331 371469
rect 154365 371409 154377 371469
rect 154319 371397 154377 371409
rect 154477 371469 154535 371481
rect 154477 371409 154489 371469
rect 154523 371409 154535 371469
rect 154477 371397 154535 371409
rect 154595 371469 154653 371481
rect 154595 371409 154607 371469
rect 154641 371409 154653 371469
rect 154595 371397 154653 371409
rect 154753 371469 154811 371481
rect 154753 371409 154765 371469
rect 154799 371409 154811 371469
rect 154753 371397 154811 371409
rect 154871 371469 154929 371481
rect 154871 371409 154883 371469
rect 154917 371409 154929 371469
rect 154871 371397 154929 371409
rect 155029 371469 155087 371481
rect 155029 371409 155041 371469
rect 155075 371409 155087 371469
rect 155029 371397 155087 371409
rect 155147 371469 155205 371481
rect 155147 371409 155159 371469
rect 155193 371409 155205 371469
rect 155147 371397 155205 371409
rect 155305 371469 155363 371481
rect 155305 371409 155317 371469
rect 155351 371409 155363 371469
rect 155305 371397 155363 371409
rect 155423 371469 155481 371481
rect 155423 371409 155435 371469
rect 155469 371409 155481 371469
rect 155423 371397 155481 371409
rect 155581 371469 155639 371481
rect 155581 371409 155593 371469
rect 155627 371409 155639 371469
rect 155581 371397 155639 371409
rect 155699 371469 155757 371481
rect 155699 371409 155711 371469
rect 155745 371409 155757 371469
rect 155699 371397 155757 371409
rect 155857 371469 155915 371481
rect 155857 371409 155869 371469
rect 155903 371409 155915 371469
rect 155857 371397 155915 371409
rect 155975 371469 156033 371481
rect 155975 371409 155987 371469
rect 156021 371409 156033 371469
rect 155975 371397 156033 371409
rect 156133 371469 156191 371481
rect 156133 371409 156145 371469
rect 156179 371409 156191 371469
rect 156133 371397 156191 371409
rect 156251 371469 156309 371481
rect 156251 371409 156263 371469
rect 156297 371409 156309 371469
rect 156251 371397 156309 371409
rect 156409 371469 156467 371481
rect 156409 371409 156421 371469
rect 156455 371409 156467 371469
rect 156409 371397 156467 371409
rect 156527 371469 156585 371481
rect 156527 371409 156539 371469
rect 156573 371409 156585 371469
rect 156527 371397 156585 371409
rect 156685 371469 156743 371481
rect 156685 371409 156697 371469
rect 156731 371409 156743 371469
rect 156685 371397 156743 371409
rect 156803 371469 156861 371481
rect 156803 371409 156815 371469
rect 156849 371409 156861 371469
rect 156803 371397 156861 371409
rect 156961 371469 157019 371481
rect 156961 371409 156973 371469
rect 157007 371409 157019 371469
rect 156961 371397 157019 371409
rect 157079 371469 157137 371481
rect 157079 371409 157091 371469
rect 157125 371409 157137 371469
rect 157079 371397 157137 371409
rect 157237 371469 157295 371481
rect 157237 371409 157249 371469
rect 157283 371409 157295 371469
rect 157237 371397 157295 371409
rect 418829 371759 418887 371771
rect 418829 371699 418841 371759
rect 418875 371699 418887 371759
rect 418829 371687 418887 371699
rect 418987 371759 419045 371771
rect 418987 371699 418999 371759
rect 419033 371699 419045 371759
rect 418987 371687 419045 371699
rect 419105 371759 419163 371771
rect 419105 371699 419117 371759
rect 419151 371699 419163 371759
rect 419105 371687 419163 371699
rect 419263 371759 419321 371771
rect 419263 371699 419275 371759
rect 419309 371699 419321 371759
rect 419263 371687 419321 371699
rect 419381 371759 419439 371771
rect 419381 371699 419393 371759
rect 419427 371699 419439 371759
rect 419381 371687 419439 371699
rect 419539 371759 419597 371771
rect 419539 371699 419551 371759
rect 419585 371699 419597 371759
rect 419539 371687 419597 371699
rect 419657 371759 419715 371771
rect 419657 371699 419669 371759
rect 419703 371699 419715 371759
rect 419657 371687 419715 371699
rect 419815 371759 419873 371771
rect 419815 371699 419827 371759
rect 419861 371699 419873 371759
rect 419815 371687 419873 371699
rect 419933 371759 419991 371771
rect 419933 371699 419945 371759
rect 419979 371699 419991 371759
rect 419933 371687 419991 371699
rect 420091 371759 420149 371771
rect 420091 371699 420103 371759
rect 420137 371699 420149 371759
rect 420091 371687 420149 371699
rect 420209 371759 420267 371771
rect 420209 371699 420221 371759
rect 420255 371699 420267 371759
rect 420209 371687 420267 371699
rect 420367 371759 420425 371771
rect 420367 371699 420379 371759
rect 420413 371699 420425 371759
rect 420367 371687 420425 371699
rect 420485 371759 420543 371771
rect 420485 371699 420497 371759
rect 420531 371699 420543 371759
rect 420485 371687 420543 371699
rect 420643 371759 420701 371771
rect 420643 371699 420655 371759
rect 420689 371699 420701 371759
rect 420643 371687 420701 371699
rect 420761 371759 420819 371771
rect 420761 371699 420773 371759
rect 420807 371699 420819 371759
rect 420761 371687 420819 371699
rect 420919 371759 420977 371771
rect 420919 371699 420931 371759
rect 420965 371699 420977 371759
rect 420919 371687 420977 371699
rect 421037 371759 421095 371771
rect 421037 371699 421049 371759
rect 421083 371699 421095 371759
rect 421037 371687 421095 371699
rect 421195 371759 421253 371771
rect 421195 371699 421207 371759
rect 421241 371699 421253 371759
rect 421195 371687 421253 371699
rect 421313 371759 421371 371771
rect 421313 371699 421325 371759
rect 421359 371699 421371 371759
rect 421313 371687 421371 371699
rect 421471 371759 421529 371771
rect 421471 371699 421483 371759
rect 421517 371699 421529 371759
rect 421471 371687 421529 371699
rect 508828 371431 508886 371443
rect 508828 371371 508840 371431
rect 508874 371371 508886 371431
rect 508828 371359 508886 371371
rect 508986 371431 509044 371443
rect 508986 371371 508998 371431
rect 509032 371371 509044 371431
rect 508986 371359 509044 371371
rect 509104 371431 509162 371443
rect 509104 371371 509116 371431
rect 509150 371371 509162 371431
rect 509104 371359 509162 371371
rect 509262 371431 509320 371443
rect 509262 371371 509274 371431
rect 509308 371371 509320 371431
rect 509262 371359 509320 371371
rect 509380 371431 509438 371443
rect 509380 371371 509392 371431
rect 509426 371371 509438 371431
rect 509380 371359 509438 371371
rect 509538 371431 509596 371443
rect 509538 371371 509550 371431
rect 509584 371371 509596 371431
rect 509538 371359 509596 371371
rect 509656 371431 509714 371443
rect 509656 371371 509668 371431
rect 509702 371371 509714 371431
rect 509656 371359 509714 371371
rect 509814 371431 509872 371443
rect 509814 371371 509826 371431
rect 509860 371371 509872 371431
rect 509814 371359 509872 371371
rect 509932 371431 509990 371443
rect 509932 371371 509944 371431
rect 509978 371371 509990 371431
rect 509932 371359 509990 371371
rect 510090 371431 510148 371443
rect 510090 371371 510102 371431
rect 510136 371371 510148 371431
rect 510090 371359 510148 371371
rect 232636 370873 232694 370885
rect 232636 370813 232648 370873
rect 232682 370813 232694 370873
rect 232636 370801 232694 370813
rect 232794 370873 232852 370885
rect 232794 370813 232806 370873
rect 232840 370813 232852 370873
rect 232794 370801 232852 370813
rect 232912 370873 232970 370885
rect 232912 370813 232924 370873
rect 232958 370813 232970 370873
rect 232912 370801 232970 370813
rect 233070 370873 233128 370885
rect 233070 370813 233082 370873
rect 233116 370813 233128 370873
rect 233070 370801 233128 370813
rect 233188 370873 233246 370885
rect 233188 370813 233200 370873
rect 233234 370813 233246 370873
rect 233188 370801 233246 370813
rect 233346 370873 233404 370885
rect 233346 370813 233358 370873
rect 233392 370813 233404 370873
rect 233346 370801 233404 370813
rect 233464 370873 233522 370885
rect 233464 370813 233476 370873
rect 233510 370813 233522 370873
rect 233464 370801 233522 370813
rect 233622 370873 233680 370885
rect 233622 370813 233634 370873
rect 233668 370813 233680 370873
rect 233622 370801 233680 370813
rect 233740 370873 233798 370885
rect 233740 370813 233752 370873
rect 233786 370813 233798 370873
rect 233740 370801 233798 370813
rect 233898 370873 233956 370885
rect 233898 370813 233910 370873
rect 233944 370813 233956 370873
rect 233898 370801 233956 370813
rect 234016 370873 234074 370885
rect 234016 370813 234028 370873
rect 234062 370813 234074 370873
rect 234016 370801 234074 370813
rect 234174 370873 234232 370885
rect 234174 370813 234186 370873
rect 234220 370813 234232 370873
rect 234174 370801 234232 370813
rect 234292 370873 234350 370885
rect 234292 370813 234304 370873
rect 234338 370813 234350 370873
rect 234292 370801 234350 370813
rect 234450 370873 234508 370885
rect 234450 370813 234462 370873
rect 234496 370813 234508 370873
rect 234450 370801 234508 370813
rect 234568 370873 234626 370885
rect 234568 370813 234580 370873
rect 234614 370813 234626 370873
rect 234568 370801 234626 370813
rect 234726 370873 234784 370885
rect 234726 370813 234738 370873
rect 234772 370813 234784 370873
rect 234726 370801 234784 370813
rect 234844 370873 234902 370885
rect 234844 370813 234856 370873
rect 234890 370813 234902 370873
rect 234844 370801 234902 370813
rect 235002 370873 235060 370885
rect 235002 370813 235014 370873
rect 235048 370813 235060 370873
rect 235002 370801 235060 370813
rect 235120 370873 235178 370885
rect 235120 370813 235132 370873
rect 235166 370813 235178 370873
rect 235120 370801 235178 370813
rect 235278 370873 235336 370885
rect 235278 370813 235290 370873
rect 235324 370813 235336 370873
rect 235278 370801 235336 370813
rect 235396 370873 235454 370885
rect 235396 370813 235408 370873
rect 235442 370813 235454 370873
rect 235396 370801 235454 370813
rect 235554 370873 235612 370885
rect 235554 370813 235566 370873
rect 235600 370813 235612 370873
rect 235554 370801 235612 370813
rect 235672 370873 235730 370885
rect 235672 370813 235684 370873
rect 235718 370813 235730 370873
rect 235672 370801 235730 370813
rect 235830 370873 235888 370885
rect 235830 370813 235842 370873
rect 235876 370813 235888 370873
rect 235830 370801 235888 370813
rect 235948 370873 236006 370885
rect 235948 370813 235960 370873
rect 235994 370813 236006 370873
rect 235948 370801 236006 370813
rect 236106 370873 236164 370885
rect 236106 370813 236118 370873
rect 236152 370813 236164 370873
rect 236106 370801 236164 370813
rect 236224 370873 236282 370885
rect 236224 370813 236236 370873
rect 236270 370813 236282 370873
rect 236224 370801 236282 370813
rect 236382 370873 236440 370885
rect 236382 370813 236394 370873
rect 236428 370813 236440 370873
rect 236382 370801 236440 370813
rect 236500 370873 236558 370885
rect 236500 370813 236512 370873
rect 236546 370813 236558 370873
rect 236500 370801 236558 370813
rect 236658 370873 236716 370885
rect 236658 370813 236670 370873
rect 236704 370813 236716 370873
rect 236658 370801 236716 370813
rect 236776 370873 236834 370885
rect 236776 370813 236788 370873
rect 236822 370813 236834 370873
rect 236776 370801 236834 370813
rect 236934 370873 236992 370885
rect 236934 370813 236946 370873
rect 236980 370813 236992 370873
rect 236934 370801 236992 370813
rect 237052 370873 237110 370885
rect 237052 370813 237064 370873
rect 237098 370813 237110 370873
rect 237052 370801 237110 370813
rect 237210 370873 237268 370885
rect 237210 370813 237222 370873
rect 237256 370813 237268 370873
rect 237210 370801 237268 370813
rect 237328 370873 237386 370885
rect 237328 370813 237340 370873
rect 237374 370813 237386 370873
rect 237328 370801 237386 370813
rect 237486 370873 237544 370885
rect 237486 370813 237498 370873
rect 237532 370813 237544 370873
rect 237486 370801 237544 370813
rect 237604 370873 237662 370885
rect 237604 370813 237616 370873
rect 237650 370813 237662 370873
rect 237604 370801 237662 370813
rect 237762 370873 237820 370885
rect 237762 370813 237774 370873
rect 237808 370813 237820 370873
rect 237762 370801 237820 370813
rect 237880 370873 237938 370885
rect 237880 370813 237892 370873
rect 237926 370813 237938 370873
rect 237880 370801 237938 370813
rect 238038 370873 238096 370885
rect 238038 370813 238050 370873
rect 238084 370813 238096 370873
rect 238038 370801 238096 370813
rect 238156 370873 238214 370885
rect 238156 370813 238168 370873
rect 238202 370813 238214 370873
rect 238156 370801 238214 370813
rect 238314 370873 238372 370885
rect 238314 370813 238326 370873
rect 238360 370813 238372 370873
rect 238314 370801 238372 370813
rect 238432 370873 238490 370885
rect 238432 370813 238444 370873
rect 238478 370813 238490 370873
rect 238432 370801 238490 370813
rect 238590 370873 238648 370885
rect 238590 370813 238602 370873
rect 238636 370813 238648 370873
rect 238590 370801 238648 370813
rect 238708 370873 238766 370885
rect 238708 370813 238720 370873
rect 238754 370813 238766 370873
rect 238708 370801 238766 370813
rect 238866 370873 238924 370885
rect 238866 370813 238878 370873
rect 238912 370813 238924 370873
rect 238866 370801 238924 370813
rect 238984 370873 239042 370885
rect 238984 370813 238996 370873
rect 239030 370813 239042 370873
rect 238984 370801 239042 370813
rect 239142 370873 239200 370885
rect 239142 370813 239154 370873
rect 239188 370813 239200 370873
rect 239142 370801 239200 370813
rect 239260 370873 239318 370885
rect 239260 370813 239272 370873
rect 239306 370813 239318 370873
rect 239260 370801 239318 370813
rect 239418 370873 239476 370885
rect 239418 370813 239430 370873
rect 239464 370813 239476 370873
rect 239418 370801 239476 370813
rect 239536 370873 239594 370885
rect 239536 370813 239548 370873
rect 239582 370813 239594 370873
rect 239536 370801 239594 370813
rect 239694 370873 239752 370885
rect 239694 370813 239706 370873
rect 239740 370813 239752 370873
rect 239694 370801 239752 370813
rect 239812 370873 239870 370885
rect 239812 370813 239824 370873
rect 239858 370813 239870 370873
rect 239812 370801 239870 370813
rect 239970 370873 240028 370885
rect 239970 370813 239982 370873
rect 240016 370813 240028 370873
rect 239970 370801 240028 370813
rect 240088 370873 240146 370885
rect 240088 370813 240100 370873
rect 240134 370813 240146 370873
rect 240088 370801 240146 370813
rect 240246 370873 240304 370885
rect 240246 370813 240258 370873
rect 240292 370813 240304 370873
rect 240246 370801 240304 370813
rect 240364 370873 240422 370885
rect 240364 370813 240376 370873
rect 240410 370813 240422 370873
rect 240364 370801 240422 370813
rect 240522 370873 240580 370885
rect 240522 370813 240534 370873
rect 240568 370813 240580 370873
rect 240522 370801 240580 370813
rect 240640 370873 240698 370885
rect 240640 370813 240652 370873
rect 240686 370813 240698 370873
rect 240640 370801 240698 370813
rect 240798 370873 240856 370885
rect 240798 370813 240810 370873
rect 240844 370813 240856 370873
rect 240798 370801 240856 370813
rect 240916 370873 240974 370885
rect 240916 370813 240928 370873
rect 240962 370813 240974 370873
rect 240916 370801 240974 370813
rect 241074 370873 241132 370885
rect 241074 370813 241086 370873
rect 241120 370813 241132 370873
rect 241074 370801 241132 370813
rect 241192 370873 241250 370885
rect 241192 370813 241204 370873
rect 241238 370813 241250 370873
rect 241192 370801 241250 370813
rect 241350 370873 241408 370885
rect 241350 370813 241362 370873
rect 241396 370813 241408 370873
rect 241350 370801 241408 370813
rect 241468 370873 241526 370885
rect 241468 370813 241480 370873
rect 241514 370813 241526 370873
rect 241468 370801 241526 370813
rect 241626 370873 241684 370885
rect 241626 370813 241638 370873
rect 241672 370813 241684 370873
rect 241626 370801 241684 370813
rect 241744 370873 241802 370885
rect 241744 370813 241756 370873
rect 241790 370813 241802 370873
rect 241744 370801 241802 370813
rect 241902 370873 241960 370885
rect 241902 370813 241914 370873
rect 241948 370813 241960 370873
rect 241902 370801 241960 370813
rect 242020 370873 242078 370885
rect 242020 370813 242032 370873
rect 242066 370813 242078 370873
rect 242020 370801 242078 370813
rect 242178 370873 242236 370885
rect 242178 370813 242190 370873
rect 242224 370813 242236 370873
rect 242178 370801 242236 370813
rect 242296 370873 242354 370885
rect 242296 370813 242308 370873
rect 242342 370813 242354 370873
rect 242296 370801 242354 370813
rect 242454 370873 242512 370885
rect 242454 370813 242466 370873
rect 242500 370813 242512 370873
rect 242454 370801 242512 370813
rect 242572 370873 242630 370885
rect 242572 370813 242584 370873
rect 242618 370813 242630 370873
rect 242572 370801 242630 370813
rect 242730 370873 242788 370885
rect 242730 370813 242742 370873
rect 242776 370813 242788 370873
rect 242730 370801 242788 370813
rect 242848 370873 242906 370885
rect 242848 370813 242860 370873
rect 242894 370813 242906 370873
rect 242848 370801 242906 370813
rect 243006 370873 243064 370885
rect 243006 370813 243018 370873
rect 243052 370813 243064 370873
rect 243006 370801 243064 370813
rect 243124 370873 243182 370885
rect 243124 370813 243136 370873
rect 243170 370813 243182 370873
rect 243124 370801 243182 370813
rect 243282 370873 243340 370885
rect 243282 370813 243294 370873
rect 243328 370813 243340 370873
rect 243282 370801 243340 370813
rect 243400 370873 243458 370885
rect 243400 370813 243412 370873
rect 243446 370813 243458 370873
rect 243400 370801 243458 370813
rect 243558 370873 243616 370885
rect 243558 370813 243570 370873
rect 243604 370813 243616 370873
rect 243558 370801 243616 370813
rect 243676 370873 243734 370885
rect 243676 370813 243688 370873
rect 243722 370813 243734 370873
rect 243676 370801 243734 370813
rect 243834 370873 243892 370885
rect 243834 370813 243846 370873
rect 243880 370813 243892 370873
rect 243834 370801 243892 370813
rect 243952 370873 244010 370885
rect 243952 370813 243964 370873
rect 243998 370813 244010 370873
rect 243952 370801 244010 370813
rect 244110 370873 244168 370885
rect 244110 370813 244122 370873
rect 244156 370813 244168 370873
rect 244110 370801 244168 370813
rect 244228 370873 244286 370885
rect 244228 370813 244240 370873
rect 244274 370813 244286 370873
rect 244228 370801 244286 370813
rect 244386 370873 244444 370885
rect 244386 370813 244398 370873
rect 244432 370813 244444 370873
rect 244386 370801 244444 370813
rect 244504 370873 244562 370885
rect 244504 370813 244516 370873
rect 244550 370813 244562 370873
rect 244504 370801 244562 370813
rect 244662 370873 244720 370885
rect 244662 370813 244674 370873
rect 244708 370813 244720 370873
rect 244662 370801 244720 370813
rect 244780 370873 244838 370885
rect 244780 370813 244792 370873
rect 244826 370813 244838 370873
rect 244780 370801 244838 370813
rect 244938 370873 244996 370885
rect 244938 370813 244950 370873
rect 244984 370813 244996 370873
rect 244938 370801 244996 370813
rect 245056 370873 245114 370885
rect 245056 370813 245068 370873
rect 245102 370813 245114 370873
rect 245056 370801 245114 370813
rect 245214 370873 245272 370885
rect 245214 370813 245226 370873
rect 245260 370813 245272 370873
rect 245214 370801 245272 370813
rect 245332 370873 245390 370885
rect 245332 370813 245344 370873
rect 245378 370813 245390 370873
rect 245332 370801 245390 370813
rect 245490 370873 245548 370885
rect 245490 370813 245502 370873
rect 245536 370813 245548 370873
rect 245490 370801 245548 370813
rect 245608 370873 245666 370885
rect 245608 370813 245620 370873
rect 245654 370813 245666 370873
rect 245608 370801 245666 370813
rect 245766 370873 245824 370885
rect 245766 370813 245778 370873
rect 245812 370813 245824 370873
rect 245766 370801 245824 370813
rect 245884 370873 245942 370885
rect 245884 370813 245896 370873
rect 245930 370813 245942 370873
rect 245884 370801 245942 370813
rect 246042 370873 246100 370885
rect 246042 370813 246054 370873
rect 246088 370813 246100 370873
rect 246042 370801 246100 370813
rect 246160 370873 246218 370885
rect 246160 370813 246172 370873
rect 246206 370813 246218 370873
rect 246160 370801 246218 370813
rect 246318 370873 246376 370885
rect 246318 370813 246330 370873
rect 246364 370813 246376 370873
rect 246318 370801 246376 370813
rect 246436 370873 246494 370885
rect 246436 370813 246448 370873
rect 246482 370813 246494 370873
rect 246436 370801 246494 370813
rect 246594 370873 246652 370885
rect 246594 370813 246606 370873
rect 246640 370813 246652 370873
rect 246594 370801 246652 370813
rect 58828 251431 58886 251443
rect 58828 251371 58840 251431
rect 58874 251371 58886 251431
rect 58828 251359 58886 251371
rect 58986 251431 59044 251443
rect 58986 251371 58998 251431
rect 59032 251371 59044 251431
rect 58986 251359 59044 251371
rect 59104 251431 59162 251443
rect 59104 251371 59116 251431
rect 59150 251371 59162 251431
rect 59104 251359 59162 251371
rect 59262 251431 59320 251443
rect 59262 251371 59274 251431
rect 59308 251371 59320 251431
rect 59262 251359 59320 251371
rect 59380 251431 59438 251443
rect 59380 251371 59392 251431
rect 59426 251371 59438 251431
rect 59380 251359 59438 251371
rect 59538 251431 59596 251443
rect 59538 251371 59550 251431
rect 59584 251371 59596 251431
rect 59538 251359 59596 251371
rect 59656 251431 59714 251443
rect 59656 251371 59668 251431
rect 59702 251371 59714 251431
rect 59656 251359 59714 251371
rect 59814 251431 59872 251443
rect 59814 251371 59826 251431
rect 59860 251371 59872 251431
rect 59814 251359 59872 251371
rect 59932 251431 59990 251443
rect 59932 251371 59944 251431
rect 59978 251371 59990 251431
rect 59932 251359 59990 251371
rect 60090 251431 60148 251443
rect 60090 251371 60102 251431
rect 60136 251371 60148 251431
rect 60090 251359 60148 251371
rect 147953 251555 148011 251567
rect 147953 251495 147965 251555
rect 147999 251495 148011 251555
rect 147953 251483 148011 251495
rect 148111 251555 148169 251567
rect 148111 251495 148123 251555
rect 148157 251495 148169 251555
rect 148111 251483 148169 251495
rect 148229 251555 148287 251567
rect 148229 251495 148241 251555
rect 148275 251495 148287 251555
rect 148229 251483 148287 251495
rect 148387 251555 148445 251567
rect 148387 251495 148399 251555
rect 148433 251495 148445 251555
rect 148387 251483 148445 251495
rect 148505 251555 148563 251567
rect 148505 251495 148517 251555
rect 148551 251495 148563 251555
rect 148505 251483 148563 251495
rect 148663 251555 148721 251567
rect 148663 251495 148675 251555
rect 148709 251495 148721 251555
rect 148663 251483 148721 251495
rect 148781 251555 148839 251567
rect 148781 251495 148793 251555
rect 148827 251495 148839 251555
rect 148781 251483 148839 251495
rect 148939 251555 148997 251567
rect 148939 251495 148951 251555
rect 148985 251495 148997 251555
rect 148939 251483 148997 251495
rect 149057 251555 149115 251567
rect 149057 251495 149069 251555
rect 149103 251495 149115 251555
rect 149057 251483 149115 251495
rect 149215 251555 149273 251567
rect 149215 251495 149227 251555
rect 149261 251495 149273 251555
rect 149215 251483 149273 251495
rect 149333 251555 149391 251567
rect 149333 251495 149345 251555
rect 149379 251495 149391 251555
rect 149333 251483 149391 251495
rect 149491 251555 149549 251567
rect 149491 251495 149503 251555
rect 149537 251495 149549 251555
rect 149491 251483 149549 251495
rect 149609 251555 149667 251567
rect 149609 251495 149621 251555
rect 149655 251495 149667 251555
rect 149609 251483 149667 251495
rect 149767 251555 149825 251567
rect 149767 251495 149779 251555
rect 149813 251495 149825 251555
rect 149767 251483 149825 251495
rect 149885 251555 149943 251567
rect 149885 251495 149897 251555
rect 149931 251495 149943 251555
rect 149885 251483 149943 251495
rect 150043 251555 150101 251567
rect 150043 251495 150055 251555
rect 150089 251495 150101 251555
rect 150043 251483 150101 251495
rect 150161 251555 150219 251567
rect 150161 251495 150173 251555
rect 150207 251495 150219 251555
rect 150161 251483 150219 251495
rect 150319 251555 150377 251567
rect 150319 251495 150331 251555
rect 150365 251495 150377 251555
rect 150319 251483 150377 251495
rect 150437 251555 150495 251567
rect 150437 251495 150449 251555
rect 150483 251495 150495 251555
rect 150437 251483 150495 251495
rect 150595 251555 150653 251567
rect 150595 251495 150607 251555
rect 150641 251495 150653 251555
rect 150595 251483 150653 251495
rect 234197 251755 234255 251767
rect 234197 251695 234209 251755
rect 234243 251695 234255 251755
rect 234197 251683 234255 251695
rect 234355 251755 234413 251767
rect 234355 251695 234367 251755
rect 234401 251695 234413 251755
rect 234355 251683 234413 251695
rect 234473 251755 234531 251767
rect 234473 251695 234485 251755
rect 234519 251695 234531 251755
rect 234473 251683 234531 251695
rect 234631 251755 234689 251767
rect 234631 251695 234643 251755
rect 234677 251695 234689 251755
rect 234631 251683 234689 251695
rect 234749 251755 234807 251767
rect 234749 251695 234761 251755
rect 234795 251695 234807 251755
rect 234749 251683 234807 251695
rect 234907 251755 234965 251767
rect 234907 251695 234919 251755
rect 234953 251695 234965 251755
rect 234907 251683 234965 251695
rect 235025 251755 235083 251767
rect 235025 251695 235037 251755
rect 235071 251695 235083 251755
rect 235025 251683 235083 251695
rect 235183 251755 235241 251767
rect 235183 251695 235195 251755
rect 235229 251695 235241 251755
rect 235183 251683 235241 251695
rect 235301 251755 235359 251767
rect 235301 251695 235313 251755
rect 235347 251695 235359 251755
rect 235301 251683 235359 251695
rect 235459 251755 235517 251767
rect 235459 251695 235471 251755
rect 235505 251695 235517 251755
rect 235459 251683 235517 251695
rect 235577 251755 235635 251767
rect 235577 251695 235589 251755
rect 235623 251695 235635 251755
rect 235577 251683 235635 251695
rect 235735 251755 235793 251767
rect 235735 251695 235747 251755
rect 235781 251695 235793 251755
rect 235735 251683 235793 251695
rect 235853 251755 235911 251767
rect 235853 251695 235865 251755
rect 235899 251695 235911 251755
rect 235853 251683 235911 251695
rect 236011 251755 236069 251767
rect 236011 251695 236023 251755
rect 236057 251695 236069 251755
rect 236011 251683 236069 251695
rect 236129 251755 236187 251767
rect 236129 251695 236141 251755
rect 236175 251695 236187 251755
rect 236129 251683 236187 251695
rect 236287 251755 236345 251767
rect 236287 251695 236299 251755
rect 236333 251695 236345 251755
rect 236287 251683 236345 251695
rect 236405 251755 236463 251767
rect 236405 251695 236417 251755
rect 236451 251695 236463 251755
rect 236405 251683 236463 251695
rect 236563 251755 236621 251767
rect 236563 251695 236575 251755
rect 236609 251695 236621 251755
rect 236563 251683 236621 251695
rect 236681 251755 236739 251767
rect 236681 251695 236693 251755
rect 236727 251695 236739 251755
rect 236681 251683 236739 251695
rect 236839 251755 236897 251767
rect 236839 251695 236851 251755
rect 236885 251695 236897 251755
rect 236839 251683 236897 251695
rect 236957 251755 237015 251767
rect 236957 251695 236969 251755
rect 237003 251695 237015 251755
rect 236957 251683 237015 251695
rect 237115 251755 237173 251767
rect 237115 251695 237127 251755
rect 237161 251695 237173 251755
rect 237115 251683 237173 251695
rect 237233 251755 237291 251767
rect 237233 251695 237245 251755
rect 237279 251695 237291 251755
rect 237233 251683 237291 251695
rect 237391 251755 237449 251767
rect 237391 251695 237403 251755
rect 237437 251695 237449 251755
rect 237391 251683 237449 251695
rect 237509 251755 237567 251767
rect 237509 251695 237521 251755
rect 237555 251695 237567 251755
rect 237509 251683 237567 251695
rect 237667 251755 237725 251767
rect 237667 251695 237679 251755
rect 237713 251695 237725 251755
rect 237667 251683 237725 251695
rect 237785 251755 237843 251767
rect 237785 251695 237797 251755
rect 237831 251695 237843 251755
rect 237785 251683 237843 251695
rect 237943 251755 238001 251767
rect 237943 251695 237955 251755
rect 237989 251695 238001 251755
rect 237943 251683 238001 251695
rect 238061 251755 238119 251767
rect 238061 251695 238073 251755
rect 238107 251695 238119 251755
rect 238061 251683 238119 251695
rect 238219 251755 238277 251767
rect 238219 251695 238231 251755
rect 238265 251695 238277 251755
rect 238219 251683 238277 251695
rect 238337 251755 238395 251767
rect 238337 251695 238349 251755
rect 238383 251695 238395 251755
rect 238337 251683 238395 251695
rect 238495 251755 238553 251767
rect 238495 251695 238507 251755
rect 238541 251695 238553 251755
rect 238495 251683 238553 251695
rect 238613 251755 238671 251767
rect 238613 251695 238625 251755
rect 238659 251695 238671 251755
rect 238613 251683 238671 251695
rect 238771 251755 238829 251767
rect 238771 251695 238783 251755
rect 238817 251695 238829 251755
rect 238771 251683 238829 251695
rect 238889 251755 238947 251767
rect 238889 251695 238901 251755
rect 238935 251695 238947 251755
rect 238889 251683 238947 251695
rect 239047 251755 239105 251767
rect 239047 251695 239059 251755
rect 239093 251695 239105 251755
rect 239047 251683 239105 251695
rect 239165 251755 239223 251767
rect 239165 251695 239177 251755
rect 239211 251695 239223 251755
rect 239165 251683 239223 251695
rect 239323 251755 239381 251767
rect 239323 251695 239335 251755
rect 239369 251695 239381 251755
rect 239323 251683 239381 251695
rect 239441 251755 239499 251767
rect 239441 251695 239453 251755
rect 239487 251695 239499 251755
rect 239441 251683 239499 251695
rect 239599 251755 239657 251767
rect 239599 251695 239611 251755
rect 239645 251695 239657 251755
rect 239599 251683 239657 251695
rect 239717 251755 239775 251767
rect 239717 251695 239729 251755
rect 239763 251695 239775 251755
rect 239717 251683 239775 251695
rect 239875 251755 239933 251767
rect 239875 251695 239887 251755
rect 239921 251695 239933 251755
rect 239875 251683 239933 251695
rect 239993 251755 240051 251767
rect 239993 251695 240005 251755
rect 240039 251695 240051 251755
rect 239993 251683 240051 251695
rect 240151 251755 240209 251767
rect 240151 251695 240163 251755
rect 240197 251695 240209 251755
rect 240151 251683 240209 251695
rect 240269 251755 240327 251767
rect 240269 251695 240281 251755
rect 240315 251695 240327 251755
rect 240269 251683 240327 251695
rect 240427 251755 240485 251767
rect 240427 251695 240439 251755
rect 240473 251695 240485 251755
rect 240427 251683 240485 251695
rect 240545 251755 240603 251767
rect 240545 251695 240557 251755
rect 240591 251695 240603 251755
rect 240545 251683 240603 251695
rect 240703 251755 240761 251767
rect 240703 251695 240715 251755
rect 240749 251695 240761 251755
rect 240703 251683 240761 251695
rect 240821 251755 240879 251767
rect 240821 251695 240833 251755
rect 240867 251695 240879 251755
rect 240821 251683 240879 251695
rect 240979 251755 241037 251767
rect 240979 251695 240991 251755
rect 241025 251695 241037 251755
rect 240979 251683 241037 251695
rect 241097 251755 241155 251767
rect 241097 251695 241109 251755
rect 241143 251695 241155 251755
rect 241097 251683 241155 251695
rect 241255 251755 241313 251767
rect 241255 251695 241267 251755
rect 241301 251695 241313 251755
rect 241255 251683 241313 251695
rect 241373 251755 241431 251767
rect 241373 251695 241385 251755
rect 241419 251695 241431 251755
rect 241373 251683 241431 251695
rect 241531 251755 241589 251767
rect 241531 251695 241543 251755
rect 241577 251695 241589 251755
rect 241531 251683 241589 251695
rect 241649 251755 241707 251767
rect 241649 251695 241661 251755
rect 241695 251695 241707 251755
rect 241649 251683 241707 251695
rect 241807 251755 241865 251767
rect 241807 251695 241819 251755
rect 241853 251695 241865 251755
rect 241807 251683 241865 251695
rect 241925 251755 241983 251767
rect 241925 251695 241937 251755
rect 241971 251695 241983 251755
rect 241925 251683 241983 251695
rect 242083 251755 242141 251767
rect 242083 251695 242095 251755
rect 242129 251695 242141 251755
rect 242083 251683 242141 251695
rect 242201 251755 242259 251767
rect 242201 251695 242213 251755
rect 242247 251695 242259 251755
rect 242201 251683 242259 251695
rect 242359 251755 242417 251767
rect 242359 251695 242371 251755
rect 242405 251695 242417 251755
rect 242359 251683 242417 251695
rect 242477 251755 242535 251767
rect 242477 251695 242489 251755
rect 242523 251695 242535 251755
rect 242477 251683 242535 251695
rect 242635 251755 242693 251767
rect 242635 251695 242647 251755
rect 242681 251695 242693 251755
rect 242635 251683 242693 251695
rect 242753 251755 242811 251767
rect 242753 251695 242765 251755
rect 242799 251695 242811 251755
rect 242753 251683 242811 251695
rect 242911 251755 242969 251767
rect 242911 251695 242923 251755
rect 242957 251695 242969 251755
rect 242911 251683 242969 251695
rect 243029 251755 243087 251767
rect 243029 251695 243041 251755
rect 243075 251695 243087 251755
rect 243029 251683 243087 251695
rect 243187 251755 243245 251767
rect 243187 251695 243199 251755
rect 243233 251695 243245 251755
rect 243187 251683 243245 251695
rect 243305 251755 243363 251767
rect 243305 251695 243317 251755
rect 243351 251695 243363 251755
rect 243305 251683 243363 251695
rect 243463 251755 243521 251767
rect 243463 251695 243475 251755
rect 243509 251695 243521 251755
rect 243463 251683 243521 251695
rect 243581 251755 243639 251767
rect 243581 251695 243593 251755
rect 243627 251695 243639 251755
rect 243581 251683 243639 251695
rect 243739 251755 243797 251767
rect 243739 251695 243751 251755
rect 243785 251695 243797 251755
rect 243739 251683 243797 251695
rect 243857 251755 243915 251767
rect 243857 251695 243869 251755
rect 243903 251695 243915 251755
rect 243857 251683 243915 251695
rect 244015 251755 244073 251767
rect 244015 251695 244027 251755
rect 244061 251695 244073 251755
rect 244015 251683 244073 251695
rect 244133 251755 244191 251767
rect 244133 251695 244145 251755
rect 244179 251695 244191 251755
rect 244133 251683 244191 251695
rect 244291 251755 244349 251767
rect 244291 251695 244303 251755
rect 244337 251695 244349 251755
rect 244291 251683 244349 251695
rect 244409 251755 244467 251767
rect 244409 251695 244421 251755
rect 244455 251695 244467 251755
rect 244409 251683 244467 251695
rect 244567 251755 244625 251767
rect 244567 251695 244579 251755
rect 244613 251695 244625 251755
rect 244567 251683 244625 251695
rect 244685 251755 244743 251767
rect 244685 251695 244697 251755
rect 244731 251695 244743 251755
rect 244685 251683 244743 251695
rect 244843 251755 244901 251767
rect 244843 251695 244855 251755
rect 244889 251695 244901 251755
rect 244843 251683 244901 251695
rect 244961 251755 245019 251767
rect 244961 251695 244973 251755
rect 245007 251695 245019 251755
rect 244961 251683 245019 251695
rect 245119 251755 245177 251767
rect 245119 251695 245131 251755
rect 245165 251695 245177 251755
rect 245119 251683 245177 251695
rect 245237 251755 245295 251767
rect 245237 251695 245249 251755
rect 245283 251695 245295 251755
rect 245237 251683 245295 251695
rect 245395 251755 245453 251767
rect 245395 251695 245407 251755
rect 245441 251695 245453 251755
rect 245395 251683 245453 251695
rect 245513 251755 245571 251767
rect 245513 251695 245525 251755
rect 245559 251695 245571 251755
rect 245513 251683 245571 251695
rect 245671 251755 245729 251767
rect 245671 251695 245683 251755
rect 245717 251695 245729 251755
rect 245671 251683 245729 251695
rect 245789 251755 245847 251767
rect 245789 251695 245801 251755
rect 245835 251695 245847 251755
rect 245789 251683 245847 251695
rect 245947 251755 246005 251767
rect 245947 251695 245959 251755
rect 245993 251695 246005 251755
rect 245947 251683 246005 251695
rect 246065 251755 246123 251767
rect 246065 251695 246077 251755
rect 246111 251695 246123 251755
rect 246065 251683 246123 251695
rect 246223 251755 246281 251767
rect 246223 251695 246235 251755
rect 246269 251695 246281 251755
rect 246223 251683 246281 251695
rect 246341 251755 246399 251767
rect 246341 251695 246353 251755
rect 246387 251695 246399 251755
rect 246341 251683 246399 251695
rect 246499 251755 246557 251767
rect 246499 251695 246511 251755
rect 246545 251695 246557 251755
rect 246499 251683 246557 251695
rect 246617 251755 246675 251767
rect 246617 251695 246629 251755
rect 246663 251695 246675 251755
rect 246617 251683 246675 251695
rect 246775 251755 246833 251767
rect 246775 251695 246787 251755
rect 246821 251695 246833 251755
rect 246775 251683 246833 251695
rect 246893 251755 246951 251767
rect 246893 251695 246905 251755
rect 246939 251695 246951 251755
rect 246893 251683 246951 251695
rect 247051 251755 247109 251767
rect 247051 251695 247063 251755
rect 247097 251695 247109 251755
rect 247051 251683 247109 251695
rect 247169 251755 247227 251767
rect 247169 251695 247181 251755
rect 247215 251695 247227 251755
rect 247169 251683 247227 251695
rect 247327 251755 247385 251767
rect 247327 251695 247339 251755
rect 247373 251695 247385 251755
rect 247327 251683 247385 251695
rect 247445 251755 247503 251767
rect 247445 251695 247457 251755
rect 247491 251695 247503 251755
rect 247445 251683 247503 251695
rect 247603 251755 247661 251767
rect 247603 251695 247615 251755
rect 247649 251695 247661 251755
rect 247603 251683 247661 251695
rect 247721 251755 247779 251767
rect 247721 251695 247733 251755
rect 247767 251695 247779 251755
rect 247721 251683 247779 251695
rect 247879 251755 247937 251767
rect 247879 251695 247891 251755
rect 247925 251695 247937 251755
rect 247879 251683 247937 251695
rect 247997 251755 248055 251767
rect 247997 251695 248009 251755
rect 248043 251695 248055 251755
rect 247997 251683 248055 251695
rect 248155 251755 248213 251767
rect 248155 251695 248167 251755
rect 248201 251695 248213 251755
rect 248155 251683 248213 251695
rect 413279 251469 413337 251481
rect 413279 251409 413291 251469
rect 413325 251409 413337 251469
rect 413279 251397 413337 251409
rect 413437 251469 413495 251481
rect 413437 251409 413449 251469
rect 413483 251409 413495 251469
rect 413437 251397 413495 251409
rect 413555 251469 413613 251481
rect 413555 251409 413567 251469
rect 413601 251409 413613 251469
rect 413555 251397 413613 251409
rect 413713 251469 413771 251481
rect 413713 251409 413725 251469
rect 413759 251409 413771 251469
rect 413713 251397 413771 251409
rect 413831 251469 413889 251481
rect 413831 251409 413843 251469
rect 413877 251409 413889 251469
rect 413831 251397 413889 251409
rect 413989 251469 414047 251481
rect 413989 251409 414001 251469
rect 414035 251409 414047 251469
rect 413989 251397 414047 251409
rect 414107 251469 414165 251481
rect 414107 251409 414119 251469
rect 414153 251409 414165 251469
rect 414107 251397 414165 251409
rect 414265 251469 414323 251481
rect 414265 251409 414277 251469
rect 414311 251409 414323 251469
rect 414265 251397 414323 251409
rect 414383 251469 414441 251481
rect 414383 251409 414395 251469
rect 414429 251409 414441 251469
rect 414383 251397 414441 251409
rect 414541 251469 414599 251481
rect 414541 251409 414553 251469
rect 414587 251409 414599 251469
rect 414541 251397 414599 251409
rect 414659 251469 414717 251481
rect 414659 251409 414671 251469
rect 414705 251409 414717 251469
rect 414659 251397 414717 251409
rect 414817 251469 414875 251481
rect 414817 251409 414829 251469
rect 414863 251409 414875 251469
rect 414817 251397 414875 251409
rect 414935 251469 414993 251481
rect 414935 251409 414947 251469
rect 414981 251409 414993 251469
rect 414935 251397 414993 251409
rect 415093 251469 415151 251481
rect 415093 251409 415105 251469
rect 415139 251409 415151 251469
rect 415093 251397 415151 251409
rect 415211 251469 415269 251481
rect 415211 251409 415223 251469
rect 415257 251409 415269 251469
rect 415211 251397 415269 251409
rect 415369 251469 415427 251481
rect 415369 251409 415381 251469
rect 415415 251409 415427 251469
rect 415369 251397 415427 251409
rect 415487 251469 415545 251481
rect 415487 251409 415499 251469
rect 415533 251409 415545 251469
rect 415487 251397 415545 251409
rect 415645 251469 415703 251481
rect 415645 251409 415657 251469
rect 415691 251409 415703 251469
rect 415645 251397 415703 251409
rect 415763 251469 415821 251481
rect 415763 251409 415775 251469
rect 415809 251409 415821 251469
rect 415763 251397 415821 251409
rect 415921 251469 415979 251481
rect 415921 251409 415933 251469
rect 415967 251409 415979 251469
rect 415921 251397 415979 251409
rect 416039 251469 416097 251481
rect 416039 251409 416051 251469
rect 416085 251409 416097 251469
rect 416039 251397 416097 251409
rect 416197 251469 416255 251481
rect 416197 251409 416209 251469
rect 416243 251409 416255 251469
rect 416197 251397 416255 251409
rect 416315 251469 416373 251481
rect 416315 251409 416327 251469
rect 416361 251409 416373 251469
rect 416315 251397 416373 251409
rect 416473 251469 416531 251481
rect 416473 251409 416485 251469
rect 416519 251409 416531 251469
rect 416473 251397 416531 251409
rect 416591 251469 416649 251481
rect 416591 251409 416603 251469
rect 416637 251409 416649 251469
rect 416591 251397 416649 251409
rect 416749 251469 416807 251481
rect 416749 251409 416761 251469
rect 416795 251409 416807 251469
rect 416749 251397 416807 251409
rect 416867 251469 416925 251481
rect 416867 251409 416879 251469
rect 416913 251409 416925 251469
rect 416867 251397 416925 251409
rect 417025 251469 417083 251481
rect 417025 251409 417037 251469
rect 417071 251409 417083 251469
rect 417025 251397 417083 251409
rect 417143 251469 417201 251481
rect 417143 251409 417155 251469
rect 417189 251409 417201 251469
rect 417143 251397 417201 251409
rect 417301 251469 417359 251481
rect 417301 251409 417313 251469
rect 417347 251409 417359 251469
rect 417301 251397 417359 251409
rect 417419 251469 417477 251481
rect 417419 251409 417431 251469
rect 417465 251409 417477 251469
rect 417419 251397 417477 251409
rect 417577 251469 417635 251481
rect 417577 251409 417589 251469
rect 417623 251409 417635 251469
rect 417577 251397 417635 251409
rect 417695 251469 417753 251481
rect 417695 251409 417707 251469
rect 417741 251409 417753 251469
rect 417695 251397 417753 251409
rect 417853 251469 417911 251481
rect 417853 251409 417865 251469
rect 417899 251409 417911 251469
rect 417853 251397 417911 251409
rect 417971 251469 418029 251481
rect 417971 251409 417983 251469
rect 418017 251409 418029 251469
rect 417971 251397 418029 251409
rect 418129 251469 418187 251481
rect 418129 251409 418141 251469
rect 418175 251409 418187 251469
rect 418129 251397 418187 251409
rect 418247 251469 418305 251481
rect 418247 251409 418259 251469
rect 418293 251409 418305 251469
rect 418247 251397 418305 251409
rect 418405 251469 418463 251481
rect 418405 251409 418417 251469
rect 418451 251409 418463 251469
rect 418405 251397 418463 251409
rect 418523 251469 418581 251481
rect 418523 251409 418535 251469
rect 418569 251409 418581 251469
rect 418523 251397 418581 251409
rect 418681 251469 418739 251481
rect 418681 251409 418693 251469
rect 418727 251409 418739 251469
rect 418681 251397 418739 251409
rect 418799 251469 418857 251481
rect 418799 251409 418811 251469
rect 418845 251409 418857 251469
rect 418799 251397 418857 251409
rect 418957 251469 419015 251481
rect 418957 251409 418969 251469
rect 419003 251409 419015 251469
rect 418957 251397 419015 251409
rect 419075 251469 419133 251481
rect 419075 251409 419087 251469
rect 419121 251409 419133 251469
rect 419075 251397 419133 251409
rect 419233 251469 419291 251481
rect 419233 251409 419245 251469
rect 419279 251409 419291 251469
rect 419233 251397 419291 251409
rect 419351 251469 419409 251481
rect 419351 251409 419363 251469
rect 419397 251409 419409 251469
rect 419351 251397 419409 251409
rect 419509 251469 419567 251481
rect 419509 251409 419521 251469
rect 419555 251409 419567 251469
rect 419509 251397 419567 251409
rect 419627 251469 419685 251481
rect 419627 251409 419639 251469
rect 419673 251409 419685 251469
rect 419627 251397 419685 251409
rect 419785 251469 419843 251481
rect 419785 251409 419797 251469
rect 419831 251409 419843 251469
rect 419785 251397 419843 251409
rect 419903 251469 419961 251481
rect 419903 251409 419915 251469
rect 419949 251409 419961 251469
rect 419903 251397 419961 251409
rect 420061 251469 420119 251481
rect 420061 251409 420073 251469
rect 420107 251409 420119 251469
rect 420061 251397 420119 251409
rect 420179 251469 420237 251481
rect 420179 251409 420191 251469
rect 420225 251409 420237 251469
rect 420179 251397 420237 251409
rect 420337 251469 420395 251481
rect 420337 251409 420349 251469
rect 420383 251409 420395 251469
rect 420337 251397 420395 251409
rect 420455 251469 420513 251481
rect 420455 251409 420467 251469
rect 420501 251409 420513 251469
rect 420455 251397 420513 251409
rect 420613 251469 420671 251481
rect 420613 251409 420625 251469
rect 420659 251409 420671 251469
rect 420613 251397 420671 251409
rect 420731 251469 420789 251481
rect 420731 251409 420743 251469
rect 420777 251409 420789 251469
rect 420731 251397 420789 251409
rect 420889 251469 420947 251481
rect 420889 251409 420901 251469
rect 420935 251409 420947 251469
rect 420889 251397 420947 251409
rect 421007 251469 421065 251481
rect 421007 251409 421019 251469
rect 421053 251409 421065 251469
rect 421007 251397 421065 251409
rect 421165 251469 421223 251481
rect 421165 251409 421177 251469
rect 421211 251409 421223 251469
rect 421165 251397 421223 251409
rect 421283 251469 421341 251481
rect 421283 251409 421295 251469
rect 421329 251409 421341 251469
rect 421283 251397 421341 251409
rect 421441 251469 421499 251481
rect 421441 251409 421453 251469
rect 421487 251409 421499 251469
rect 421441 251397 421499 251409
rect 421559 251469 421617 251481
rect 421559 251409 421571 251469
rect 421605 251409 421617 251469
rect 421559 251397 421617 251409
rect 421717 251469 421775 251481
rect 421717 251409 421729 251469
rect 421763 251409 421775 251469
rect 421717 251397 421775 251409
rect 421835 251469 421893 251481
rect 421835 251409 421847 251469
rect 421881 251409 421893 251469
rect 421835 251397 421893 251409
rect 421993 251469 422051 251481
rect 421993 251409 422005 251469
rect 422039 251409 422051 251469
rect 421993 251397 422051 251409
rect 422111 251469 422169 251481
rect 422111 251409 422123 251469
rect 422157 251409 422169 251469
rect 422111 251397 422169 251409
rect 422269 251469 422327 251481
rect 422269 251409 422281 251469
rect 422315 251409 422327 251469
rect 422269 251397 422327 251409
rect 422387 251469 422445 251481
rect 422387 251409 422399 251469
rect 422433 251409 422445 251469
rect 422387 251397 422445 251409
rect 422545 251469 422603 251481
rect 422545 251409 422557 251469
rect 422591 251409 422603 251469
rect 422545 251397 422603 251409
rect 422663 251469 422721 251481
rect 422663 251409 422675 251469
rect 422709 251409 422721 251469
rect 422663 251397 422721 251409
rect 422821 251469 422879 251481
rect 422821 251409 422833 251469
rect 422867 251409 422879 251469
rect 422821 251397 422879 251409
rect 422939 251469 422997 251481
rect 422939 251409 422951 251469
rect 422985 251409 422997 251469
rect 422939 251397 422997 251409
rect 423097 251469 423155 251481
rect 423097 251409 423109 251469
rect 423143 251409 423155 251469
rect 423097 251397 423155 251409
rect 423215 251469 423273 251481
rect 423215 251409 423227 251469
rect 423261 251409 423273 251469
rect 423215 251397 423273 251409
rect 423373 251469 423431 251481
rect 423373 251409 423385 251469
rect 423419 251409 423431 251469
rect 423373 251397 423431 251409
rect 423491 251469 423549 251481
rect 423491 251409 423503 251469
rect 423537 251409 423549 251469
rect 423491 251397 423549 251409
rect 423649 251469 423707 251481
rect 423649 251409 423661 251469
rect 423695 251409 423707 251469
rect 423649 251397 423707 251409
rect 423767 251469 423825 251481
rect 423767 251409 423779 251469
rect 423813 251409 423825 251469
rect 423767 251397 423825 251409
rect 423925 251469 423983 251481
rect 423925 251409 423937 251469
rect 423971 251409 423983 251469
rect 423925 251397 423983 251409
rect 424043 251469 424101 251481
rect 424043 251409 424055 251469
rect 424089 251409 424101 251469
rect 424043 251397 424101 251409
rect 424201 251469 424259 251481
rect 424201 251409 424213 251469
rect 424247 251409 424259 251469
rect 424201 251397 424259 251409
rect 424319 251469 424377 251481
rect 424319 251409 424331 251469
rect 424365 251409 424377 251469
rect 424319 251397 424377 251409
rect 424477 251469 424535 251481
rect 424477 251409 424489 251469
rect 424523 251409 424535 251469
rect 424477 251397 424535 251409
rect 424595 251469 424653 251481
rect 424595 251409 424607 251469
rect 424641 251409 424653 251469
rect 424595 251397 424653 251409
rect 424753 251469 424811 251481
rect 424753 251409 424765 251469
rect 424799 251409 424811 251469
rect 424753 251397 424811 251409
rect 424871 251469 424929 251481
rect 424871 251409 424883 251469
rect 424917 251409 424929 251469
rect 424871 251397 424929 251409
rect 425029 251469 425087 251481
rect 425029 251409 425041 251469
rect 425075 251409 425087 251469
rect 425029 251397 425087 251409
rect 425147 251469 425205 251481
rect 425147 251409 425159 251469
rect 425193 251409 425205 251469
rect 425147 251397 425205 251409
rect 425305 251469 425363 251481
rect 425305 251409 425317 251469
rect 425351 251409 425363 251469
rect 425305 251397 425363 251409
rect 425423 251469 425481 251481
rect 425423 251409 425435 251469
rect 425469 251409 425481 251469
rect 425423 251397 425481 251409
rect 425581 251469 425639 251481
rect 425581 251409 425593 251469
rect 425627 251409 425639 251469
rect 425581 251397 425639 251409
rect 425699 251469 425757 251481
rect 425699 251409 425711 251469
rect 425745 251409 425757 251469
rect 425699 251397 425757 251409
rect 425857 251469 425915 251481
rect 425857 251409 425869 251469
rect 425903 251409 425915 251469
rect 425857 251397 425915 251409
rect 425975 251469 426033 251481
rect 425975 251409 425987 251469
rect 426021 251409 426033 251469
rect 425975 251397 426033 251409
rect 426133 251469 426191 251481
rect 426133 251409 426145 251469
rect 426179 251409 426191 251469
rect 426133 251397 426191 251409
rect 426251 251469 426309 251481
rect 426251 251409 426263 251469
rect 426297 251409 426309 251469
rect 426251 251397 426309 251409
rect 426409 251469 426467 251481
rect 426409 251409 426421 251469
rect 426455 251409 426467 251469
rect 426409 251397 426467 251409
rect 426527 251469 426585 251481
rect 426527 251409 426539 251469
rect 426573 251409 426585 251469
rect 426527 251397 426585 251409
rect 426685 251469 426743 251481
rect 426685 251409 426697 251469
rect 426731 251409 426743 251469
rect 426685 251397 426743 251409
rect 426803 251469 426861 251481
rect 426803 251409 426815 251469
rect 426849 251409 426861 251469
rect 426803 251397 426861 251409
rect 426961 251469 427019 251481
rect 426961 251409 426973 251469
rect 427007 251409 427019 251469
rect 426961 251397 427019 251409
rect 427079 251469 427137 251481
rect 427079 251409 427091 251469
rect 427125 251409 427137 251469
rect 427079 251397 427137 251409
rect 427237 251469 427295 251481
rect 427237 251409 427249 251469
rect 427283 251409 427295 251469
rect 427237 251397 427295 251409
rect 503279 251469 503337 251481
rect 503279 251409 503291 251469
rect 503325 251409 503337 251469
rect 503279 251397 503337 251409
rect 503437 251469 503495 251481
rect 503437 251409 503449 251469
rect 503483 251409 503495 251469
rect 503437 251397 503495 251409
rect 503555 251469 503613 251481
rect 503555 251409 503567 251469
rect 503601 251409 503613 251469
rect 503555 251397 503613 251409
rect 503713 251469 503771 251481
rect 503713 251409 503725 251469
rect 503759 251409 503771 251469
rect 503713 251397 503771 251409
rect 503831 251469 503889 251481
rect 503831 251409 503843 251469
rect 503877 251409 503889 251469
rect 503831 251397 503889 251409
rect 503989 251469 504047 251481
rect 503989 251409 504001 251469
rect 504035 251409 504047 251469
rect 503989 251397 504047 251409
rect 504107 251469 504165 251481
rect 504107 251409 504119 251469
rect 504153 251409 504165 251469
rect 504107 251397 504165 251409
rect 504265 251469 504323 251481
rect 504265 251409 504277 251469
rect 504311 251409 504323 251469
rect 504265 251397 504323 251409
rect 504383 251469 504441 251481
rect 504383 251409 504395 251469
rect 504429 251409 504441 251469
rect 504383 251397 504441 251409
rect 504541 251469 504599 251481
rect 504541 251409 504553 251469
rect 504587 251409 504599 251469
rect 504541 251397 504599 251409
rect 504659 251469 504717 251481
rect 504659 251409 504671 251469
rect 504705 251409 504717 251469
rect 504659 251397 504717 251409
rect 504817 251469 504875 251481
rect 504817 251409 504829 251469
rect 504863 251409 504875 251469
rect 504817 251397 504875 251409
rect 504935 251469 504993 251481
rect 504935 251409 504947 251469
rect 504981 251409 504993 251469
rect 504935 251397 504993 251409
rect 505093 251469 505151 251481
rect 505093 251409 505105 251469
rect 505139 251409 505151 251469
rect 505093 251397 505151 251409
rect 505211 251469 505269 251481
rect 505211 251409 505223 251469
rect 505257 251409 505269 251469
rect 505211 251397 505269 251409
rect 505369 251469 505427 251481
rect 505369 251409 505381 251469
rect 505415 251409 505427 251469
rect 505369 251397 505427 251409
rect 505487 251469 505545 251481
rect 505487 251409 505499 251469
rect 505533 251409 505545 251469
rect 505487 251397 505545 251409
rect 505645 251469 505703 251481
rect 505645 251409 505657 251469
rect 505691 251409 505703 251469
rect 505645 251397 505703 251409
rect 505763 251469 505821 251481
rect 505763 251409 505775 251469
rect 505809 251409 505821 251469
rect 505763 251397 505821 251409
rect 505921 251469 505979 251481
rect 505921 251409 505933 251469
rect 505967 251409 505979 251469
rect 505921 251397 505979 251409
rect 506039 251469 506097 251481
rect 506039 251409 506051 251469
rect 506085 251409 506097 251469
rect 506039 251397 506097 251409
rect 506197 251469 506255 251481
rect 506197 251409 506209 251469
rect 506243 251409 506255 251469
rect 506197 251397 506255 251409
rect 506315 251469 506373 251481
rect 506315 251409 506327 251469
rect 506361 251409 506373 251469
rect 506315 251397 506373 251409
rect 506473 251469 506531 251481
rect 506473 251409 506485 251469
rect 506519 251409 506531 251469
rect 506473 251397 506531 251409
rect 506591 251469 506649 251481
rect 506591 251409 506603 251469
rect 506637 251409 506649 251469
rect 506591 251397 506649 251409
rect 506749 251469 506807 251481
rect 506749 251409 506761 251469
rect 506795 251409 506807 251469
rect 506749 251397 506807 251409
rect 506867 251469 506925 251481
rect 506867 251409 506879 251469
rect 506913 251409 506925 251469
rect 506867 251397 506925 251409
rect 507025 251469 507083 251481
rect 507025 251409 507037 251469
rect 507071 251409 507083 251469
rect 507025 251397 507083 251409
rect 507143 251469 507201 251481
rect 507143 251409 507155 251469
rect 507189 251409 507201 251469
rect 507143 251397 507201 251409
rect 507301 251469 507359 251481
rect 507301 251409 507313 251469
rect 507347 251409 507359 251469
rect 507301 251397 507359 251409
rect 507419 251469 507477 251481
rect 507419 251409 507431 251469
rect 507465 251409 507477 251469
rect 507419 251397 507477 251409
rect 507577 251469 507635 251481
rect 507577 251409 507589 251469
rect 507623 251409 507635 251469
rect 507577 251397 507635 251409
rect 507695 251469 507753 251481
rect 507695 251409 507707 251469
rect 507741 251409 507753 251469
rect 507695 251397 507753 251409
rect 507853 251469 507911 251481
rect 507853 251409 507865 251469
rect 507899 251409 507911 251469
rect 507853 251397 507911 251409
rect 507971 251469 508029 251481
rect 507971 251409 507983 251469
rect 508017 251409 508029 251469
rect 507971 251397 508029 251409
rect 508129 251469 508187 251481
rect 508129 251409 508141 251469
rect 508175 251409 508187 251469
rect 508129 251397 508187 251409
rect 508247 251469 508305 251481
rect 508247 251409 508259 251469
rect 508293 251409 508305 251469
rect 508247 251397 508305 251409
rect 508405 251469 508463 251481
rect 508405 251409 508417 251469
rect 508451 251409 508463 251469
rect 508405 251397 508463 251409
rect 508523 251469 508581 251481
rect 508523 251409 508535 251469
rect 508569 251409 508581 251469
rect 508523 251397 508581 251409
rect 508681 251469 508739 251481
rect 508681 251409 508693 251469
rect 508727 251409 508739 251469
rect 508681 251397 508739 251409
rect 508799 251469 508857 251481
rect 508799 251409 508811 251469
rect 508845 251409 508857 251469
rect 508799 251397 508857 251409
rect 508957 251469 509015 251481
rect 508957 251409 508969 251469
rect 509003 251409 509015 251469
rect 508957 251397 509015 251409
rect 509075 251469 509133 251481
rect 509075 251409 509087 251469
rect 509121 251409 509133 251469
rect 509075 251397 509133 251409
rect 509233 251469 509291 251481
rect 509233 251409 509245 251469
rect 509279 251409 509291 251469
rect 509233 251397 509291 251409
rect 509351 251469 509409 251481
rect 509351 251409 509363 251469
rect 509397 251409 509409 251469
rect 509351 251397 509409 251409
rect 509509 251469 509567 251481
rect 509509 251409 509521 251469
rect 509555 251409 509567 251469
rect 509509 251397 509567 251409
rect 509627 251469 509685 251481
rect 509627 251409 509639 251469
rect 509673 251409 509685 251469
rect 509627 251397 509685 251409
rect 509785 251469 509843 251481
rect 509785 251409 509797 251469
rect 509831 251409 509843 251469
rect 509785 251397 509843 251409
rect 509903 251469 509961 251481
rect 509903 251409 509915 251469
rect 509949 251409 509961 251469
rect 509903 251397 509961 251409
rect 510061 251469 510119 251481
rect 510061 251409 510073 251469
rect 510107 251409 510119 251469
rect 510061 251397 510119 251409
rect 510179 251469 510237 251481
rect 510179 251409 510191 251469
rect 510225 251409 510237 251469
rect 510179 251397 510237 251409
rect 510337 251469 510395 251481
rect 510337 251409 510349 251469
rect 510383 251409 510395 251469
rect 510337 251397 510395 251409
rect 510455 251469 510513 251481
rect 510455 251409 510467 251469
rect 510501 251409 510513 251469
rect 510455 251397 510513 251409
rect 510613 251469 510671 251481
rect 510613 251409 510625 251469
rect 510659 251409 510671 251469
rect 510613 251397 510671 251409
rect 510731 251469 510789 251481
rect 510731 251409 510743 251469
rect 510777 251409 510789 251469
rect 510731 251397 510789 251409
rect 510889 251469 510947 251481
rect 510889 251409 510901 251469
rect 510935 251409 510947 251469
rect 510889 251397 510947 251409
rect 511007 251469 511065 251481
rect 511007 251409 511019 251469
rect 511053 251409 511065 251469
rect 511007 251397 511065 251409
rect 511165 251469 511223 251481
rect 511165 251409 511177 251469
rect 511211 251409 511223 251469
rect 511165 251397 511223 251409
rect 511283 251469 511341 251481
rect 511283 251409 511295 251469
rect 511329 251409 511341 251469
rect 511283 251397 511341 251409
rect 511441 251469 511499 251481
rect 511441 251409 511453 251469
rect 511487 251409 511499 251469
rect 511441 251397 511499 251409
rect 511559 251469 511617 251481
rect 511559 251409 511571 251469
rect 511605 251409 511617 251469
rect 511559 251397 511617 251409
rect 511717 251469 511775 251481
rect 511717 251409 511729 251469
rect 511763 251409 511775 251469
rect 511717 251397 511775 251409
rect 511835 251469 511893 251481
rect 511835 251409 511847 251469
rect 511881 251409 511893 251469
rect 511835 251397 511893 251409
rect 511993 251469 512051 251481
rect 511993 251409 512005 251469
rect 512039 251409 512051 251469
rect 511993 251397 512051 251409
rect 512111 251469 512169 251481
rect 512111 251409 512123 251469
rect 512157 251409 512169 251469
rect 512111 251397 512169 251409
rect 512269 251469 512327 251481
rect 512269 251409 512281 251469
rect 512315 251409 512327 251469
rect 512269 251397 512327 251409
rect 512387 251469 512445 251481
rect 512387 251409 512399 251469
rect 512433 251409 512445 251469
rect 512387 251397 512445 251409
rect 512545 251469 512603 251481
rect 512545 251409 512557 251469
rect 512591 251409 512603 251469
rect 512545 251397 512603 251409
rect 512663 251469 512721 251481
rect 512663 251409 512675 251469
rect 512709 251409 512721 251469
rect 512663 251397 512721 251409
rect 512821 251469 512879 251481
rect 512821 251409 512833 251469
rect 512867 251409 512879 251469
rect 512821 251397 512879 251409
rect 512939 251469 512997 251481
rect 512939 251409 512951 251469
rect 512985 251409 512997 251469
rect 512939 251397 512997 251409
rect 513097 251469 513155 251481
rect 513097 251409 513109 251469
rect 513143 251409 513155 251469
rect 513097 251397 513155 251409
rect 513215 251469 513273 251481
rect 513215 251409 513227 251469
rect 513261 251409 513273 251469
rect 513215 251397 513273 251409
rect 513373 251469 513431 251481
rect 513373 251409 513385 251469
rect 513419 251409 513431 251469
rect 513373 251397 513431 251409
rect 513491 251469 513549 251481
rect 513491 251409 513503 251469
rect 513537 251409 513549 251469
rect 513491 251397 513549 251409
rect 513649 251469 513707 251481
rect 513649 251409 513661 251469
rect 513695 251409 513707 251469
rect 513649 251397 513707 251409
rect 513767 251469 513825 251481
rect 513767 251409 513779 251469
rect 513813 251409 513825 251469
rect 513767 251397 513825 251409
rect 513925 251469 513983 251481
rect 513925 251409 513937 251469
rect 513971 251409 513983 251469
rect 513925 251397 513983 251409
rect 514043 251469 514101 251481
rect 514043 251409 514055 251469
rect 514089 251409 514101 251469
rect 514043 251397 514101 251409
rect 514201 251469 514259 251481
rect 514201 251409 514213 251469
rect 514247 251409 514259 251469
rect 514201 251397 514259 251409
rect 514319 251469 514377 251481
rect 514319 251409 514331 251469
rect 514365 251409 514377 251469
rect 514319 251397 514377 251409
rect 514477 251469 514535 251481
rect 514477 251409 514489 251469
rect 514523 251409 514535 251469
rect 514477 251397 514535 251409
rect 514595 251469 514653 251481
rect 514595 251409 514607 251469
rect 514641 251409 514653 251469
rect 514595 251397 514653 251409
rect 514753 251469 514811 251481
rect 514753 251409 514765 251469
rect 514799 251409 514811 251469
rect 514753 251397 514811 251409
rect 514871 251469 514929 251481
rect 514871 251409 514883 251469
rect 514917 251409 514929 251469
rect 514871 251397 514929 251409
rect 515029 251469 515087 251481
rect 515029 251409 515041 251469
rect 515075 251409 515087 251469
rect 515029 251397 515087 251409
rect 515147 251469 515205 251481
rect 515147 251409 515159 251469
rect 515193 251409 515205 251469
rect 515147 251397 515205 251409
rect 515305 251469 515363 251481
rect 515305 251409 515317 251469
rect 515351 251409 515363 251469
rect 515305 251397 515363 251409
rect 515423 251469 515481 251481
rect 515423 251409 515435 251469
rect 515469 251409 515481 251469
rect 515423 251397 515481 251409
rect 515581 251469 515639 251481
rect 515581 251409 515593 251469
rect 515627 251409 515639 251469
rect 515581 251397 515639 251409
rect 515699 251469 515757 251481
rect 515699 251409 515711 251469
rect 515745 251409 515757 251469
rect 515699 251397 515757 251409
rect 515857 251469 515915 251481
rect 515857 251409 515869 251469
rect 515903 251409 515915 251469
rect 515857 251397 515915 251409
rect 515975 251469 516033 251481
rect 515975 251409 515987 251469
rect 516021 251409 516033 251469
rect 515975 251397 516033 251409
rect 516133 251469 516191 251481
rect 516133 251409 516145 251469
rect 516179 251409 516191 251469
rect 516133 251397 516191 251409
rect 516251 251469 516309 251481
rect 516251 251409 516263 251469
rect 516297 251409 516309 251469
rect 516251 251397 516309 251409
rect 516409 251469 516467 251481
rect 516409 251409 516421 251469
rect 516455 251409 516467 251469
rect 516409 251397 516467 251409
rect 516527 251469 516585 251481
rect 516527 251409 516539 251469
rect 516573 251409 516585 251469
rect 516527 251397 516585 251409
rect 516685 251469 516743 251481
rect 516685 251409 516697 251469
rect 516731 251409 516743 251469
rect 516685 251397 516743 251409
rect 516803 251469 516861 251481
rect 516803 251409 516815 251469
rect 516849 251409 516861 251469
rect 516803 251397 516861 251409
rect 516961 251469 517019 251481
rect 516961 251409 516973 251469
rect 517007 251409 517019 251469
rect 516961 251397 517019 251409
rect 517079 251469 517137 251481
rect 517079 251409 517091 251469
rect 517125 251409 517137 251469
rect 517079 251397 517137 251409
rect 517237 251469 517295 251481
rect 517237 251409 517249 251469
rect 517283 251409 517295 251469
rect 517237 251397 517295 251409
rect 322636 250873 322694 250885
rect 322636 250813 322648 250873
rect 322682 250813 322694 250873
rect 322636 250801 322694 250813
rect 322794 250873 322852 250885
rect 322794 250813 322806 250873
rect 322840 250813 322852 250873
rect 322794 250801 322852 250813
rect 322912 250873 322970 250885
rect 322912 250813 322924 250873
rect 322958 250813 322970 250873
rect 322912 250801 322970 250813
rect 323070 250873 323128 250885
rect 323070 250813 323082 250873
rect 323116 250813 323128 250873
rect 323070 250801 323128 250813
rect 323188 250873 323246 250885
rect 323188 250813 323200 250873
rect 323234 250813 323246 250873
rect 323188 250801 323246 250813
rect 323346 250873 323404 250885
rect 323346 250813 323358 250873
rect 323392 250813 323404 250873
rect 323346 250801 323404 250813
rect 323464 250873 323522 250885
rect 323464 250813 323476 250873
rect 323510 250813 323522 250873
rect 323464 250801 323522 250813
rect 323622 250873 323680 250885
rect 323622 250813 323634 250873
rect 323668 250813 323680 250873
rect 323622 250801 323680 250813
rect 323740 250873 323798 250885
rect 323740 250813 323752 250873
rect 323786 250813 323798 250873
rect 323740 250801 323798 250813
rect 323898 250873 323956 250885
rect 323898 250813 323910 250873
rect 323944 250813 323956 250873
rect 323898 250801 323956 250813
rect 324016 250873 324074 250885
rect 324016 250813 324028 250873
rect 324062 250813 324074 250873
rect 324016 250801 324074 250813
rect 324174 250873 324232 250885
rect 324174 250813 324186 250873
rect 324220 250813 324232 250873
rect 324174 250801 324232 250813
rect 324292 250873 324350 250885
rect 324292 250813 324304 250873
rect 324338 250813 324350 250873
rect 324292 250801 324350 250813
rect 324450 250873 324508 250885
rect 324450 250813 324462 250873
rect 324496 250813 324508 250873
rect 324450 250801 324508 250813
rect 324568 250873 324626 250885
rect 324568 250813 324580 250873
rect 324614 250813 324626 250873
rect 324568 250801 324626 250813
rect 324726 250873 324784 250885
rect 324726 250813 324738 250873
rect 324772 250813 324784 250873
rect 324726 250801 324784 250813
rect 324844 250873 324902 250885
rect 324844 250813 324856 250873
rect 324890 250813 324902 250873
rect 324844 250801 324902 250813
rect 325002 250873 325060 250885
rect 325002 250813 325014 250873
rect 325048 250813 325060 250873
rect 325002 250801 325060 250813
rect 325120 250873 325178 250885
rect 325120 250813 325132 250873
rect 325166 250813 325178 250873
rect 325120 250801 325178 250813
rect 325278 250873 325336 250885
rect 325278 250813 325290 250873
rect 325324 250813 325336 250873
rect 325278 250801 325336 250813
rect 325396 250873 325454 250885
rect 325396 250813 325408 250873
rect 325442 250813 325454 250873
rect 325396 250801 325454 250813
rect 325554 250873 325612 250885
rect 325554 250813 325566 250873
rect 325600 250813 325612 250873
rect 325554 250801 325612 250813
rect 325672 250873 325730 250885
rect 325672 250813 325684 250873
rect 325718 250813 325730 250873
rect 325672 250801 325730 250813
rect 325830 250873 325888 250885
rect 325830 250813 325842 250873
rect 325876 250813 325888 250873
rect 325830 250801 325888 250813
rect 325948 250873 326006 250885
rect 325948 250813 325960 250873
rect 325994 250813 326006 250873
rect 325948 250801 326006 250813
rect 326106 250873 326164 250885
rect 326106 250813 326118 250873
rect 326152 250813 326164 250873
rect 326106 250801 326164 250813
rect 326224 250873 326282 250885
rect 326224 250813 326236 250873
rect 326270 250813 326282 250873
rect 326224 250801 326282 250813
rect 326382 250873 326440 250885
rect 326382 250813 326394 250873
rect 326428 250813 326440 250873
rect 326382 250801 326440 250813
rect 326500 250873 326558 250885
rect 326500 250813 326512 250873
rect 326546 250813 326558 250873
rect 326500 250801 326558 250813
rect 326658 250873 326716 250885
rect 326658 250813 326670 250873
rect 326704 250813 326716 250873
rect 326658 250801 326716 250813
rect 326776 250873 326834 250885
rect 326776 250813 326788 250873
rect 326822 250813 326834 250873
rect 326776 250801 326834 250813
rect 326934 250873 326992 250885
rect 326934 250813 326946 250873
rect 326980 250813 326992 250873
rect 326934 250801 326992 250813
rect 327052 250873 327110 250885
rect 327052 250813 327064 250873
rect 327098 250813 327110 250873
rect 327052 250801 327110 250813
rect 327210 250873 327268 250885
rect 327210 250813 327222 250873
rect 327256 250813 327268 250873
rect 327210 250801 327268 250813
rect 327328 250873 327386 250885
rect 327328 250813 327340 250873
rect 327374 250813 327386 250873
rect 327328 250801 327386 250813
rect 327486 250873 327544 250885
rect 327486 250813 327498 250873
rect 327532 250813 327544 250873
rect 327486 250801 327544 250813
rect 327604 250873 327662 250885
rect 327604 250813 327616 250873
rect 327650 250813 327662 250873
rect 327604 250801 327662 250813
rect 327762 250873 327820 250885
rect 327762 250813 327774 250873
rect 327808 250813 327820 250873
rect 327762 250801 327820 250813
rect 327880 250873 327938 250885
rect 327880 250813 327892 250873
rect 327926 250813 327938 250873
rect 327880 250801 327938 250813
rect 328038 250873 328096 250885
rect 328038 250813 328050 250873
rect 328084 250813 328096 250873
rect 328038 250801 328096 250813
rect 328156 250873 328214 250885
rect 328156 250813 328168 250873
rect 328202 250813 328214 250873
rect 328156 250801 328214 250813
rect 328314 250873 328372 250885
rect 328314 250813 328326 250873
rect 328360 250813 328372 250873
rect 328314 250801 328372 250813
rect 328432 250873 328490 250885
rect 328432 250813 328444 250873
rect 328478 250813 328490 250873
rect 328432 250801 328490 250813
rect 328590 250873 328648 250885
rect 328590 250813 328602 250873
rect 328636 250813 328648 250873
rect 328590 250801 328648 250813
rect 328708 250873 328766 250885
rect 328708 250813 328720 250873
rect 328754 250813 328766 250873
rect 328708 250801 328766 250813
rect 328866 250873 328924 250885
rect 328866 250813 328878 250873
rect 328912 250813 328924 250873
rect 328866 250801 328924 250813
rect 328984 250873 329042 250885
rect 328984 250813 328996 250873
rect 329030 250813 329042 250873
rect 328984 250801 329042 250813
rect 329142 250873 329200 250885
rect 329142 250813 329154 250873
rect 329188 250813 329200 250873
rect 329142 250801 329200 250813
rect 329260 250873 329318 250885
rect 329260 250813 329272 250873
rect 329306 250813 329318 250873
rect 329260 250801 329318 250813
rect 329418 250873 329476 250885
rect 329418 250813 329430 250873
rect 329464 250813 329476 250873
rect 329418 250801 329476 250813
rect 329536 250873 329594 250885
rect 329536 250813 329548 250873
rect 329582 250813 329594 250873
rect 329536 250801 329594 250813
rect 329694 250873 329752 250885
rect 329694 250813 329706 250873
rect 329740 250813 329752 250873
rect 329694 250801 329752 250813
rect 329812 250873 329870 250885
rect 329812 250813 329824 250873
rect 329858 250813 329870 250873
rect 329812 250801 329870 250813
rect 329970 250873 330028 250885
rect 329970 250813 329982 250873
rect 330016 250813 330028 250873
rect 329970 250801 330028 250813
rect 330088 250873 330146 250885
rect 330088 250813 330100 250873
rect 330134 250813 330146 250873
rect 330088 250801 330146 250813
rect 330246 250873 330304 250885
rect 330246 250813 330258 250873
rect 330292 250813 330304 250873
rect 330246 250801 330304 250813
rect 330364 250873 330422 250885
rect 330364 250813 330376 250873
rect 330410 250813 330422 250873
rect 330364 250801 330422 250813
rect 330522 250873 330580 250885
rect 330522 250813 330534 250873
rect 330568 250813 330580 250873
rect 330522 250801 330580 250813
rect 330640 250873 330698 250885
rect 330640 250813 330652 250873
rect 330686 250813 330698 250873
rect 330640 250801 330698 250813
rect 330798 250873 330856 250885
rect 330798 250813 330810 250873
rect 330844 250813 330856 250873
rect 330798 250801 330856 250813
rect 330916 250873 330974 250885
rect 330916 250813 330928 250873
rect 330962 250813 330974 250873
rect 330916 250801 330974 250813
rect 331074 250873 331132 250885
rect 331074 250813 331086 250873
rect 331120 250813 331132 250873
rect 331074 250801 331132 250813
rect 331192 250873 331250 250885
rect 331192 250813 331204 250873
rect 331238 250813 331250 250873
rect 331192 250801 331250 250813
rect 331350 250873 331408 250885
rect 331350 250813 331362 250873
rect 331396 250813 331408 250873
rect 331350 250801 331408 250813
rect 331468 250873 331526 250885
rect 331468 250813 331480 250873
rect 331514 250813 331526 250873
rect 331468 250801 331526 250813
rect 331626 250873 331684 250885
rect 331626 250813 331638 250873
rect 331672 250813 331684 250873
rect 331626 250801 331684 250813
rect 331744 250873 331802 250885
rect 331744 250813 331756 250873
rect 331790 250813 331802 250873
rect 331744 250801 331802 250813
rect 331902 250873 331960 250885
rect 331902 250813 331914 250873
rect 331948 250813 331960 250873
rect 331902 250801 331960 250813
rect 332020 250873 332078 250885
rect 332020 250813 332032 250873
rect 332066 250813 332078 250873
rect 332020 250801 332078 250813
rect 332178 250873 332236 250885
rect 332178 250813 332190 250873
rect 332224 250813 332236 250873
rect 332178 250801 332236 250813
rect 332296 250873 332354 250885
rect 332296 250813 332308 250873
rect 332342 250813 332354 250873
rect 332296 250801 332354 250813
rect 332454 250873 332512 250885
rect 332454 250813 332466 250873
rect 332500 250813 332512 250873
rect 332454 250801 332512 250813
rect 332572 250873 332630 250885
rect 332572 250813 332584 250873
rect 332618 250813 332630 250873
rect 332572 250801 332630 250813
rect 332730 250873 332788 250885
rect 332730 250813 332742 250873
rect 332776 250813 332788 250873
rect 332730 250801 332788 250813
rect 332848 250873 332906 250885
rect 332848 250813 332860 250873
rect 332894 250813 332906 250873
rect 332848 250801 332906 250813
rect 333006 250873 333064 250885
rect 333006 250813 333018 250873
rect 333052 250813 333064 250873
rect 333006 250801 333064 250813
rect 333124 250873 333182 250885
rect 333124 250813 333136 250873
rect 333170 250813 333182 250873
rect 333124 250801 333182 250813
rect 333282 250873 333340 250885
rect 333282 250813 333294 250873
rect 333328 250813 333340 250873
rect 333282 250801 333340 250813
rect 333400 250873 333458 250885
rect 333400 250813 333412 250873
rect 333446 250813 333458 250873
rect 333400 250801 333458 250813
rect 333558 250873 333616 250885
rect 333558 250813 333570 250873
rect 333604 250813 333616 250873
rect 333558 250801 333616 250813
rect 333676 250873 333734 250885
rect 333676 250813 333688 250873
rect 333722 250813 333734 250873
rect 333676 250801 333734 250813
rect 333834 250873 333892 250885
rect 333834 250813 333846 250873
rect 333880 250813 333892 250873
rect 333834 250801 333892 250813
rect 333952 250873 334010 250885
rect 333952 250813 333964 250873
rect 333998 250813 334010 250873
rect 333952 250801 334010 250813
rect 334110 250873 334168 250885
rect 334110 250813 334122 250873
rect 334156 250813 334168 250873
rect 334110 250801 334168 250813
rect 334228 250873 334286 250885
rect 334228 250813 334240 250873
rect 334274 250813 334286 250873
rect 334228 250801 334286 250813
rect 334386 250873 334444 250885
rect 334386 250813 334398 250873
rect 334432 250813 334444 250873
rect 334386 250801 334444 250813
rect 334504 250873 334562 250885
rect 334504 250813 334516 250873
rect 334550 250813 334562 250873
rect 334504 250801 334562 250813
rect 334662 250873 334720 250885
rect 334662 250813 334674 250873
rect 334708 250813 334720 250873
rect 334662 250801 334720 250813
rect 334780 250873 334838 250885
rect 334780 250813 334792 250873
rect 334826 250813 334838 250873
rect 334780 250801 334838 250813
rect 334938 250873 334996 250885
rect 334938 250813 334950 250873
rect 334984 250813 334996 250873
rect 334938 250801 334996 250813
rect 335056 250873 335114 250885
rect 335056 250813 335068 250873
rect 335102 250813 335114 250873
rect 335056 250801 335114 250813
rect 335214 250873 335272 250885
rect 335214 250813 335226 250873
rect 335260 250813 335272 250873
rect 335214 250801 335272 250813
rect 335332 250873 335390 250885
rect 335332 250813 335344 250873
rect 335378 250813 335390 250873
rect 335332 250801 335390 250813
rect 335490 250873 335548 250885
rect 335490 250813 335502 250873
rect 335536 250813 335548 250873
rect 335490 250801 335548 250813
rect 335608 250873 335666 250885
rect 335608 250813 335620 250873
rect 335654 250813 335666 250873
rect 335608 250801 335666 250813
rect 335766 250873 335824 250885
rect 335766 250813 335778 250873
rect 335812 250813 335824 250873
rect 335766 250801 335824 250813
rect 335884 250873 335942 250885
rect 335884 250813 335896 250873
rect 335930 250813 335942 250873
rect 335884 250801 335942 250813
rect 336042 250873 336100 250885
rect 336042 250813 336054 250873
rect 336088 250813 336100 250873
rect 336042 250801 336100 250813
rect 336160 250873 336218 250885
rect 336160 250813 336172 250873
rect 336206 250813 336218 250873
rect 336160 250801 336218 250813
rect 336318 250873 336376 250885
rect 336318 250813 336330 250873
rect 336364 250813 336376 250873
rect 336318 250801 336376 250813
rect 336436 250873 336494 250885
rect 336436 250813 336448 250873
rect 336482 250813 336494 250873
rect 336436 250801 336494 250813
rect 336594 250873 336652 250885
rect 336594 250813 336606 250873
rect 336640 250813 336652 250873
rect 336594 250801 336652 250813
rect 149553 55971 149611 55983
rect 149553 55795 149565 55971
rect 149599 55795 149611 55971
rect 149553 55783 149611 55795
rect 149711 55971 149769 55983
rect 149711 55795 149723 55971
rect 149757 55795 149769 55971
rect 149711 55783 149769 55795
rect 239563 55681 239621 55693
rect 239563 55505 239575 55681
rect 239609 55505 239621 55681
rect 239563 55493 239621 55505
rect 239721 55681 239779 55693
rect 239721 55505 239733 55681
rect 239767 55505 239779 55681
rect 239721 55493 239779 55505
rect 419553 55971 419611 55983
rect 419553 55795 419565 55971
rect 419599 55795 419611 55971
rect 419553 55783 419611 55795
rect 419711 55971 419769 55983
rect 419711 55795 419723 55971
rect 419757 55795 419769 55971
rect 419711 55783 419769 55795
rect 509563 55681 509621 55693
rect 509563 55505 509575 55681
rect 509609 55505 509621 55681
rect 509563 55493 509621 55505
rect 509721 55681 509779 55693
rect 509721 55505 509733 55681
rect 509767 55505 509779 55681
rect 509721 55493 509779 55505
<< mvpdiff >>
rect 419265 657454 419323 657466
rect 419265 657278 419277 657454
rect 419311 657278 419323 657454
rect 419265 657266 419323 657278
rect 419423 657454 419481 657466
rect 419423 657278 419435 657454
rect 419469 657278 419481 657454
rect 419423 657266 419481 657278
rect 329463 580530 329521 580542
rect 329463 580354 329475 580530
rect 329509 580354 329521 580530
rect 329463 580342 329521 580354
rect 329621 580530 329679 580542
rect 329621 580354 329633 580530
rect 329667 580354 329679 580530
rect 329621 580342 329679 580354
rect 149463 145530 149521 145542
rect 149463 145354 149475 145530
rect 149509 145354 149521 145530
rect 149463 145342 149521 145354
rect 149621 145530 149679 145542
rect 149621 145354 149633 145530
rect 149667 145354 149679 145530
rect 149621 145342 149679 145354
rect 419463 145530 419521 145542
rect 419463 145354 419475 145530
rect 419509 145354 419521 145530
rect 419463 145342 419521 145354
rect 419621 145530 419679 145542
rect 419621 145354 419633 145530
rect 419667 145354 419679 145530
rect 419621 145342 419679 145354
<< ndiffc >>
rect 329114 657720 329148 657896
rect 329202 657720 329236 657896
rect 509114 657720 509148 657896
rect 509202 657720 509236 657896
rect 149312 655796 149346 655972
rect 149400 655796 149434 655972
rect 239312 580796 239346 580972
rect 239400 580796 239434 580972
rect 239312 145796 239346 145972
rect 239400 145796 239434 145972
rect 509312 145796 509346 145972
rect 509400 145796 509434 145972
rect 59312 55796 59346 55972
rect 59400 55796 59434 55972
rect 329312 55796 329346 55972
rect 329400 55796 329434 55972
<< pdiffc >>
rect 239295 655758 239329 655934
rect 239383 655758 239417 655934
rect 59295 145758 59329 145934
rect 59383 145758 59417 145934
rect 329295 145758 329329 145934
rect 329383 145758 329417 145934
<< mvndiffc >>
rect 59565 655795 59599 655971
rect 59723 655795 59757 655971
rect 419367 582719 419401 582895
rect 419525 582719 419559 582895
rect 509377 582429 509411 582605
rect 509535 582429 509569 582605
rect 59565 580795 59599 580971
rect 59723 580795 59757 580971
rect 149575 580505 149609 580681
rect 149733 580505 149767 580681
rect 58841 491699 58875 491759
rect 58999 491699 59033 491759
rect 59117 491699 59151 491759
rect 59275 491699 59309 491759
rect 59393 491699 59427 491759
rect 59551 491699 59585 491759
rect 59669 491699 59703 491759
rect 59827 491699 59861 491759
rect 59945 491699 59979 491759
rect 60103 491699 60137 491759
rect 60221 491699 60255 491759
rect 60379 491699 60413 491759
rect 60497 491699 60531 491759
rect 60655 491699 60689 491759
rect 60773 491699 60807 491759
rect 60931 491699 60965 491759
rect 61049 491699 61083 491759
rect 61207 491699 61241 491759
rect 61325 491699 61359 491759
rect 61483 491699 61517 491759
rect 323831 492087 323865 492147
rect 323989 492087 324023 492147
rect 324107 492087 324141 492147
rect 324265 492087 324299 492147
rect 324383 492087 324417 492147
rect 324541 492087 324575 492147
rect 324659 492087 324693 492147
rect 324817 492087 324851 492147
rect 324935 492087 324969 492147
rect 325093 492087 325127 492147
rect 325211 492087 325245 492147
rect 325369 492087 325403 492147
rect 325487 492087 325521 492147
rect 325645 492087 325679 492147
rect 325763 492087 325797 492147
rect 325921 492087 325955 492147
rect 326039 492087 326073 492147
rect 326197 492087 326231 492147
rect 326315 492087 326349 492147
rect 326473 492087 326507 492147
rect 326591 492087 326625 492147
rect 326749 492087 326783 492147
rect 326867 492087 326901 492147
rect 327025 492087 327059 492147
rect 327143 492087 327177 492147
rect 327301 492087 327335 492147
rect 327419 492087 327453 492147
rect 327577 492087 327611 492147
rect 327695 492087 327729 492147
rect 327853 492087 327887 492147
rect 327971 492087 328005 492147
rect 328129 492087 328163 492147
rect 328247 492087 328281 492147
rect 328405 492087 328439 492147
rect 328523 492087 328557 492147
rect 328681 492087 328715 492147
rect 328799 492087 328833 492147
rect 328957 492087 328991 492147
rect 329075 492087 329109 492147
rect 329233 492087 329267 492147
rect 329351 492087 329385 492147
rect 329509 492087 329543 492147
rect 329627 492087 329661 492147
rect 329785 492087 329819 492147
rect 329903 492087 329937 492147
rect 330061 492087 330095 492147
rect 330179 492087 330213 492147
rect 330337 492087 330371 492147
rect 330455 492087 330489 492147
rect 330613 492087 330647 492147
rect 330731 492087 330765 492147
rect 330889 492087 330923 492147
rect 331007 492087 331041 492147
rect 331165 492087 331199 492147
rect 331283 492087 331317 492147
rect 331441 492087 331475 492147
rect 331559 492087 331593 492147
rect 331717 492087 331751 492147
rect 331835 492087 331869 492147
rect 331993 492087 332027 492147
rect 332111 492087 332145 492147
rect 332269 492087 332303 492147
rect 332387 492087 332421 492147
rect 332545 492087 332579 492147
rect 332663 492087 332697 492147
rect 332821 492087 332855 492147
rect 332939 492087 332973 492147
rect 333097 492087 333131 492147
rect 333215 492087 333249 492147
rect 333373 492087 333407 492147
rect 333491 492087 333525 492147
rect 333649 492087 333683 492147
rect 333767 492087 333801 492147
rect 333925 492087 333959 492147
rect 334043 492087 334077 492147
rect 334201 492087 334235 492147
rect 334319 492087 334353 492147
rect 334477 492087 334511 492147
rect 334595 492087 334629 492147
rect 334753 492087 334787 492147
rect 334871 492087 334905 492147
rect 335029 492087 335063 492147
rect 335147 492087 335181 492147
rect 335305 492087 335339 492147
rect 335423 492087 335457 492147
rect 335581 492087 335615 492147
rect 335699 492087 335733 492147
rect 335857 492087 335891 492147
rect 335975 492087 336009 492147
rect 336133 492087 336167 492147
rect 336251 492087 336285 492147
rect 336409 492087 336443 492147
rect 336527 492087 336561 492147
rect 336685 492087 336719 492147
rect 336803 492087 336837 492147
rect 336961 492087 336995 492147
rect 337079 492087 337113 492147
rect 337237 492087 337271 492147
rect 337355 492087 337389 492147
rect 337513 492087 337547 492147
rect 337631 492087 337665 492147
rect 337789 492087 337823 492147
rect 143291 491409 143325 491469
rect 143449 491409 143483 491469
rect 143567 491409 143601 491469
rect 143725 491409 143759 491469
rect 143843 491409 143877 491469
rect 144001 491409 144035 491469
rect 144119 491409 144153 491469
rect 144277 491409 144311 491469
rect 144395 491409 144429 491469
rect 144553 491409 144587 491469
rect 144671 491409 144705 491469
rect 144829 491409 144863 491469
rect 144947 491409 144981 491469
rect 145105 491409 145139 491469
rect 145223 491409 145257 491469
rect 145381 491409 145415 491469
rect 145499 491409 145533 491469
rect 145657 491409 145691 491469
rect 145775 491409 145809 491469
rect 145933 491409 145967 491469
rect 146051 491409 146085 491469
rect 146209 491409 146243 491469
rect 146327 491409 146361 491469
rect 146485 491409 146519 491469
rect 146603 491409 146637 491469
rect 146761 491409 146795 491469
rect 146879 491409 146913 491469
rect 147037 491409 147071 491469
rect 147155 491409 147189 491469
rect 147313 491409 147347 491469
rect 147431 491409 147465 491469
rect 147589 491409 147623 491469
rect 147707 491409 147741 491469
rect 147865 491409 147899 491469
rect 147983 491409 148017 491469
rect 148141 491409 148175 491469
rect 148259 491409 148293 491469
rect 148417 491409 148451 491469
rect 148535 491409 148569 491469
rect 148693 491409 148727 491469
rect 148811 491409 148845 491469
rect 148969 491409 149003 491469
rect 149087 491409 149121 491469
rect 149245 491409 149279 491469
rect 149363 491409 149397 491469
rect 149521 491409 149555 491469
rect 149639 491409 149673 491469
rect 149797 491409 149831 491469
rect 149915 491409 149949 491469
rect 150073 491409 150107 491469
rect 150191 491409 150225 491469
rect 150349 491409 150383 491469
rect 150467 491409 150501 491469
rect 150625 491409 150659 491469
rect 150743 491409 150777 491469
rect 150901 491409 150935 491469
rect 151019 491409 151053 491469
rect 151177 491409 151211 491469
rect 151295 491409 151329 491469
rect 151453 491409 151487 491469
rect 151571 491409 151605 491469
rect 151729 491409 151763 491469
rect 151847 491409 151881 491469
rect 152005 491409 152039 491469
rect 152123 491409 152157 491469
rect 152281 491409 152315 491469
rect 152399 491409 152433 491469
rect 152557 491409 152591 491469
rect 152675 491409 152709 491469
rect 152833 491409 152867 491469
rect 152951 491409 152985 491469
rect 153109 491409 153143 491469
rect 153227 491409 153261 491469
rect 153385 491409 153419 491469
rect 153503 491409 153537 491469
rect 153661 491409 153695 491469
rect 153779 491409 153813 491469
rect 153937 491409 153971 491469
rect 154055 491409 154089 491469
rect 154213 491409 154247 491469
rect 154331 491409 154365 491469
rect 154489 491409 154523 491469
rect 154607 491409 154641 491469
rect 154765 491409 154799 491469
rect 154883 491409 154917 491469
rect 155041 491409 155075 491469
rect 155159 491409 155193 491469
rect 155317 491409 155351 491469
rect 155435 491409 155469 491469
rect 155593 491409 155627 491469
rect 155711 491409 155745 491469
rect 155869 491409 155903 491469
rect 155987 491409 156021 491469
rect 156145 491409 156179 491469
rect 156263 491409 156297 491469
rect 156421 491409 156455 491469
rect 156539 491409 156573 491469
rect 156697 491409 156731 491469
rect 156815 491409 156849 491469
rect 156973 491409 157007 491469
rect 157091 491409 157125 491469
rect 157249 491409 157283 491469
rect 418840 491371 418874 491431
rect 418998 491371 419032 491431
rect 419116 491371 419150 491431
rect 419274 491371 419308 491431
rect 419392 491371 419426 491431
rect 419550 491371 419584 491431
rect 419668 491371 419702 491431
rect 419826 491371 419860 491431
rect 419944 491371 419978 491431
rect 420102 491371 420136 491431
rect 508841 491699 508875 491759
rect 508999 491699 509033 491759
rect 509117 491699 509151 491759
rect 509275 491699 509309 491759
rect 509393 491699 509427 491759
rect 509551 491699 509585 491759
rect 509669 491699 509703 491759
rect 509827 491699 509861 491759
rect 509945 491699 509979 491759
rect 510103 491699 510137 491759
rect 510221 491699 510255 491759
rect 510379 491699 510413 491759
rect 510497 491699 510531 491759
rect 510655 491699 510689 491759
rect 510773 491699 510807 491759
rect 510931 491699 510965 491759
rect 511049 491699 511083 491759
rect 511207 491699 511241 491759
rect 511325 491699 511359 491759
rect 511483 491699 511517 491759
rect 232648 490813 232682 490873
rect 232806 490813 232840 490873
rect 232924 490813 232958 490873
rect 233082 490813 233116 490873
rect 233200 490813 233234 490873
rect 233358 490813 233392 490873
rect 233476 490813 233510 490873
rect 233634 490813 233668 490873
rect 233752 490813 233786 490873
rect 233910 490813 233944 490873
rect 234028 490813 234062 490873
rect 234186 490813 234220 490873
rect 234304 490813 234338 490873
rect 234462 490813 234496 490873
rect 234580 490813 234614 490873
rect 234738 490813 234772 490873
rect 234856 490813 234890 490873
rect 235014 490813 235048 490873
rect 235132 490813 235166 490873
rect 235290 490813 235324 490873
rect 235408 490813 235442 490873
rect 235566 490813 235600 490873
rect 235684 490813 235718 490873
rect 235842 490813 235876 490873
rect 235960 490813 235994 490873
rect 236118 490813 236152 490873
rect 236236 490813 236270 490873
rect 236394 490813 236428 490873
rect 236512 490813 236546 490873
rect 236670 490813 236704 490873
rect 236788 490813 236822 490873
rect 236946 490813 236980 490873
rect 237064 490813 237098 490873
rect 237222 490813 237256 490873
rect 237340 490813 237374 490873
rect 237498 490813 237532 490873
rect 237616 490813 237650 490873
rect 237774 490813 237808 490873
rect 237892 490813 237926 490873
rect 238050 490813 238084 490873
rect 238168 490813 238202 490873
rect 238326 490813 238360 490873
rect 238444 490813 238478 490873
rect 238602 490813 238636 490873
rect 238720 490813 238754 490873
rect 238878 490813 238912 490873
rect 238996 490813 239030 490873
rect 239154 490813 239188 490873
rect 239272 490813 239306 490873
rect 239430 490813 239464 490873
rect 239548 490813 239582 490873
rect 239706 490813 239740 490873
rect 239824 490813 239858 490873
rect 239982 490813 240016 490873
rect 240100 490813 240134 490873
rect 240258 490813 240292 490873
rect 240376 490813 240410 490873
rect 240534 490813 240568 490873
rect 240652 490813 240686 490873
rect 240810 490813 240844 490873
rect 240928 490813 240962 490873
rect 241086 490813 241120 490873
rect 241204 490813 241238 490873
rect 241362 490813 241396 490873
rect 241480 490813 241514 490873
rect 241638 490813 241672 490873
rect 241756 490813 241790 490873
rect 241914 490813 241948 490873
rect 242032 490813 242066 490873
rect 242190 490813 242224 490873
rect 242308 490813 242342 490873
rect 242466 490813 242500 490873
rect 242584 490813 242618 490873
rect 242742 490813 242776 490873
rect 242860 490813 242894 490873
rect 243018 490813 243052 490873
rect 243136 490813 243170 490873
rect 243294 490813 243328 490873
rect 243412 490813 243446 490873
rect 243570 490813 243604 490873
rect 243688 490813 243722 490873
rect 243846 490813 243880 490873
rect 243964 490813 243998 490873
rect 244122 490813 244156 490873
rect 244240 490813 244274 490873
rect 244398 490813 244432 490873
rect 244516 490813 244550 490873
rect 244674 490813 244708 490873
rect 244792 490813 244826 490873
rect 244950 490813 244984 490873
rect 245068 490813 245102 490873
rect 245226 490813 245260 490873
rect 245344 490813 245378 490873
rect 245502 490813 245536 490873
rect 245620 490813 245654 490873
rect 245778 490813 245812 490873
rect 245896 490813 245930 490873
rect 246054 490813 246088 490873
rect 246172 490813 246206 490873
rect 246330 490813 246364 490873
rect 246448 490813 246482 490873
rect 246606 490813 246640 490873
rect 323831 372087 323865 372147
rect 323989 372087 324023 372147
rect 324107 372087 324141 372147
rect 324265 372087 324299 372147
rect 324383 372087 324417 372147
rect 324541 372087 324575 372147
rect 324659 372087 324693 372147
rect 324817 372087 324851 372147
rect 324935 372087 324969 372147
rect 325093 372087 325127 372147
rect 325211 372087 325245 372147
rect 325369 372087 325403 372147
rect 325487 372087 325521 372147
rect 325645 372087 325679 372147
rect 325763 372087 325797 372147
rect 325921 372087 325955 372147
rect 326039 372087 326073 372147
rect 326197 372087 326231 372147
rect 326315 372087 326349 372147
rect 326473 372087 326507 372147
rect 326591 372087 326625 372147
rect 326749 372087 326783 372147
rect 326867 372087 326901 372147
rect 327025 372087 327059 372147
rect 327143 372087 327177 372147
rect 327301 372087 327335 372147
rect 327419 372087 327453 372147
rect 327577 372087 327611 372147
rect 327695 372087 327729 372147
rect 327853 372087 327887 372147
rect 327971 372087 328005 372147
rect 328129 372087 328163 372147
rect 328247 372087 328281 372147
rect 328405 372087 328439 372147
rect 328523 372087 328557 372147
rect 328681 372087 328715 372147
rect 328799 372087 328833 372147
rect 328957 372087 328991 372147
rect 329075 372087 329109 372147
rect 329233 372087 329267 372147
rect 329351 372087 329385 372147
rect 329509 372087 329543 372147
rect 329627 372087 329661 372147
rect 329785 372087 329819 372147
rect 329903 372087 329937 372147
rect 330061 372087 330095 372147
rect 330179 372087 330213 372147
rect 330337 372087 330371 372147
rect 330455 372087 330489 372147
rect 330613 372087 330647 372147
rect 330731 372087 330765 372147
rect 330889 372087 330923 372147
rect 331007 372087 331041 372147
rect 331165 372087 331199 372147
rect 331283 372087 331317 372147
rect 331441 372087 331475 372147
rect 331559 372087 331593 372147
rect 331717 372087 331751 372147
rect 331835 372087 331869 372147
rect 331993 372087 332027 372147
rect 332111 372087 332145 372147
rect 332269 372087 332303 372147
rect 332387 372087 332421 372147
rect 332545 372087 332579 372147
rect 332663 372087 332697 372147
rect 332821 372087 332855 372147
rect 332939 372087 332973 372147
rect 333097 372087 333131 372147
rect 333215 372087 333249 372147
rect 333373 372087 333407 372147
rect 333491 372087 333525 372147
rect 333649 372087 333683 372147
rect 333767 372087 333801 372147
rect 333925 372087 333959 372147
rect 334043 372087 334077 372147
rect 334201 372087 334235 372147
rect 334319 372087 334353 372147
rect 334477 372087 334511 372147
rect 334595 372087 334629 372147
rect 334753 372087 334787 372147
rect 334871 372087 334905 372147
rect 335029 372087 335063 372147
rect 335147 372087 335181 372147
rect 335305 372087 335339 372147
rect 335423 372087 335457 372147
rect 335581 372087 335615 372147
rect 335699 372087 335733 372147
rect 335857 372087 335891 372147
rect 335975 372087 336009 372147
rect 336133 372087 336167 372147
rect 336251 372087 336285 372147
rect 336409 372087 336443 372147
rect 336527 372087 336561 372147
rect 336685 372087 336719 372147
rect 336803 372087 336837 372147
rect 336961 372087 336995 372147
rect 337079 372087 337113 372147
rect 337237 372087 337271 372147
rect 337355 372087 337389 372147
rect 337513 372087 337547 372147
rect 337631 372087 337665 372147
rect 337789 372087 337823 372147
rect 53291 371409 53325 371469
rect 53449 371409 53483 371469
rect 53567 371409 53601 371469
rect 53725 371409 53759 371469
rect 53843 371409 53877 371469
rect 54001 371409 54035 371469
rect 54119 371409 54153 371469
rect 54277 371409 54311 371469
rect 54395 371409 54429 371469
rect 54553 371409 54587 371469
rect 54671 371409 54705 371469
rect 54829 371409 54863 371469
rect 54947 371409 54981 371469
rect 55105 371409 55139 371469
rect 55223 371409 55257 371469
rect 55381 371409 55415 371469
rect 55499 371409 55533 371469
rect 55657 371409 55691 371469
rect 55775 371409 55809 371469
rect 55933 371409 55967 371469
rect 56051 371409 56085 371469
rect 56209 371409 56243 371469
rect 56327 371409 56361 371469
rect 56485 371409 56519 371469
rect 56603 371409 56637 371469
rect 56761 371409 56795 371469
rect 56879 371409 56913 371469
rect 57037 371409 57071 371469
rect 57155 371409 57189 371469
rect 57313 371409 57347 371469
rect 57431 371409 57465 371469
rect 57589 371409 57623 371469
rect 57707 371409 57741 371469
rect 57865 371409 57899 371469
rect 57983 371409 58017 371469
rect 58141 371409 58175 371469
rect 58259 371409 58293 371469
rect 58417 371409 58451 371469
rect 58535 371409 58569 371469
rect 58693 371409 58727 371469
rect 58811 371409 58845 371469
rect 58969 371409 59003 371469
rect 59087 371409 59121 371469
rect 59245 371409 59279 371469
rect 59363 371409 59397 371469
rect 59521 371409 59555 371469
rect 59639 371409 59673 371469
rect 59797 371409 59831 371469
rect 59915 371409 59949 371469
rect 60073 371409 60107 371469
rect 60191 371409 60225 371469
rect 60349 371409 60383 371469
rect 60467 371409 60501 371469
rect 60625 371409 60659 371469
rect 60743 371409 60777 371469
rect 60901 371409 60935 371469
rect 61019 371409 61053 371469
rect 61177 371409 61211 371469
rect 61295 371409 61329 371469
rect 61453 371409 61487 371469
rect 61571 371409 61605 371469
rect 61729 371409 61763 371469
rect 61847 371409 61881 371469
rect 62005 371409 62039 371469
rect 62123 371409 62157 371469
rect 62281 371409 62315 371469
rect 62399 371409 62433 371469
rect 62557 371409 62591 371469
rect 62675 371409 62709 371469
rect 62833 371409 62867 371469
rect 62951 371409 62985 371469
rect 63109 371409 63143 371469
rect 63227 371409 63261 371469
rect 63385 371409 63419 371469
rect 63503 371409 63537 371469
rect 63661 371409 63695 371469
rect 63779 371409 63813 371469
rect 63937 371409 63971 371469
rect 64055 371409 64089 371469
rect 64213 371409 64247 371469
rect 64331 371409 64365 371469
rect 64489 371409 64523 371469
rect 64607 371409 64641 371469
rect 64765 371409 64799 371469
rect 64883 371409 64917 371469
rect 65041 371409 65075 371469
rect 65159 371409 65193 371469
rect 65317 371409 65351 371469
rect 65435 371409 65469 371469
rect 65593 371409 65627 371469
rect 65711 371409 65745 371469
rect 65869 371409 65903 371469
rect 65987 371409 66021 371469
rect 66145 371409 66179 371469
rect 66263 371409 66297 371469
rect 66421 371409 66455 371469
rect 66539 371409 66573 371469
rect 66697 371409 66731 371469
rect 66815 371409 66849 371469
rect 66973 371409 67007 371469
rect 67091 371409 67125 371469
rect 67249 371409 67283 371469
rect 143291 371409 143325 371469
rect 143449 371409 143483 371469
rect 143567 371409 143601 371469
rect 143725 371409 143759 371469
rect 143843 371409 143877 371469
rect 144001 371409 144035 371469
rect 144119 371409 144153 371469
rect 144277 371409 144311 371469
rect 144395 371409 144429 371469
rect 144553 371409 144587 371469
rect 144671 371409 144705 371469
rect 144829 371409 144863 371469
rect 144947 371409 144981 371469
rect 145105 371409 145139 371469
rect 145223 371409 145257 371469
rect 145381 371409 145415 371469
rect 145499 371409 145533 371469
rect 145657 371409 145691 371469
rect 145775 371409 145809 371469
rect 145933 371409 145967 371469
rect 146051 371409 146085 371469
rect 146209 371409 146243 371469
rect 146327 371409 146361 371469
rect 146485 371409 146519 371469
rect 146603 371409 146637 371469
rect 146761 371409 146795 371469
rect 146879 371409 146913 371469
rect 147037 371409 147071 371469
rect 147155 371409 147189 371469
rect 147313 371409 147347 371469
rect 147431 371409 147465 371469
rect 147589 371409 147623 371469
rect 147707 371409 147741 371469
rect 147865 371409 147899 371469
rect 147983 371409 148017 371469
rect 148141 371409 148175 371469
rect 148259 371409 148293 371469
rect 148417 371409 148451 371469
rect 148535 371409 148569 371469
rect 148693 371409 148727 371469
rect 148811 371409 148845 371469
rect 148969 371409 149003 371469
rect 149087 371409 149121 371469
rect 149245 371409 149279 371469
rect 149363 371409 149397 371469
rect 149521 371409 149555 371469
rect 149639 371409 149673 371469
rect 149797 371409 149831 371469
rect 149915 371409 149949 371469
rect 150073 371409 150107 371469
rect 150191 371409 150225 371469
rect 150349 371409 150383 371469
rect 150467 371409 150501 371469
rect 150625 371409 150659 371469
rect 150743 371409 150777 371469
rect 150901 371409 150935 371469
rect 151019 371409 151053 371469
rect 151177 371409 151211 371469
rect 151295 371409 151329 371469
rect 151453 371409 151487 371469
rect 151571 371409 151605 371469
rect 151729 371409 151763 371469
rect 151847 371409 151881 371469
rect 152005 371409 152039 371469
rect 152123 371409 152157 371469
rect 152281 371409 152315 371469
rect 152399 371409 152433 371469
rect 152557 371409 152591 371469
rect 152675 371409 152709 371469
rect 152833 371409 152867 371469
rect 152951 371409 152985 371469
rect 153109 371409 153143 371469
rect 153227 371409 153261 371469
rect 153385 371409 153419 371469
rect 153503 371409 153537 371469
rect 153661 371409 153695 371469
rect 153779 371409 153813 371469
rect 153937 371409 153971 371469
rect 154055 371409 154089 371469
rect 154213 371409 154247 371469
rect 154331 371409 154365 371469
rect 154489 371409 154523 371469
rect 154607 371409 154641 371469
rect 154765 371409 154799 371469
rect 154883 371409 154917 371469
rect 155041 371409 155075 371469
rect 155159 371409 155193 371469
rect 155317 371409 155351 371469
rect 155435 371409 155469 371469
rect 155593 371409 155627 371469
rect 155711 371409 155745 371469
rect 155869 371409 155903 371469
rect 155987 371409 156021 371469
rect 156145 371409 156179 371469
rect 156263 371409 156297 371469
rect 156421 371409 156455 371469
rect 156539 371409 156573 371469
rect 156697 371409 156731 371469
rect 156815 371409 156849 371469
rect 156973 371409 157007 371469
rect 157091 371409 157125 371469
rect 157249 371409 157283 371469
rect 418841 371699 418875 371759
rect 418999 371699 419033 371759
rect 419117 371699 419151 371759
rect 419275 371699 419309 371759
rect 419393 371699 419427 371759
rect 419551 371699 419585 371759
rect 419669 371699 419703 371759
rect 419827 371699 419861 371759
rect 419945 371699 419979 371759
rect 420103 371699 420137 371759
rect 420221 371699 420255 371759
rect 420379 371699 420413 371759
rect 420497 371699 420531 371759
rect 420655 371699 420689 371759
rect 420773 371699 420807 371759
rect 420931 371699 420965 371759
rect 421049 371699 421083 371759
rect 421207 371699 421241 371759
rect 421325 371699 421359 371759
rect 421483 371699 421517 371759
rect 508840 371371 508874 371431
rect 508998 371371 509032 371431
rect 509116 371371 509150 371431
rect 509274 371371 509308 371431
rect 509392 371371 509426 371431
rect 509550 371371 509584 371431
rect 509668 371371 509702 371431
rect 509826 371371 509860 371431
rect 509944 371371 509978 371431
rect 510102 371371 510136 371431
rect 232648 370813 232682 370873
rect 232806 370813 232840 370873
rect 232924 370813 232958 370873
rect 233082 370813 233116 370873
rect 233200 370813 233234 370873
rect 233358 370813 233392 370873
rect 233476 370813 233510 370873
rect 233634 370813 233668 370873
rect 233752 370813 233786 370873
rect 233910 370813 233944 370873
rect 234028 370813 234062 370873
rect 234186 370813 234220 370873
rect 234304 370813 234338 370873
rect 234462 370813 234496 370873
rect 234580 370813 234614 370873
rect 234738 370813 234772 370873
rect 234856 370813 234890 370873
rect 235014 370813 235048 370873
rect 235132 370813 235166 370873
rect 235290 370813 235324 370873
rect 235408 370813 235442 370873
rect 235566 370813 235600 370873
rect 235684 370813 235718 370873
rect 235842 370813 235876 370873
rect 235960 370813 235994 370873
rect 236118 370813 236152 370873
rect 236236 370813 236270 370873
rect 236394 370813 236428 370873
rect 236512 370813 236546 370873
rect 236670 370813 236704 370873
rect 236788 370813 236822 370873
rect 236946 370813 236980 370873
rect 237064 370813 237098 370873
rect 237222 370813 237256 370873
rect 237340 370813 237374 370873
rect 237498 370813 237532 370873
rect 237616 370813 237650 370873
rect 237774 370813 237808 370873
rect 237892 370813 237926 370873
rect 238050 370813 238084 370873
rect 238168 370813 238202 370873
rect 238326 370813 238360 370873
rect 238444 370813 238478 370873
rect 238602 370813 238636 370873
rect 238720 370813 238754 370873
rect 238878 370813 238912 370873
rect 238996 370813 239030 370873
rect 239154 370813 239188 370873
rect 239272 370813 239306 370873
rect 239430 370813 239464 370873
rect 239548 370813 239582 370873
rect 239706 370813 239740 370873
rect 239824 370813 239858 370873
rect 239982 370813 240016 370873
rect 240100 370813 240134 370873
rect 240258 370813 240292 370873
rect 240376 370813 240410 370873
rect 240534 370813 240568 370873
rect 240652 370813 240686 370873
rect 240810 370813 240844 370873
rect 240928 370813 240962 370873
rect 241086 370813 241120 370873
rect 241204 370813 241238 370873
rect 241362 370813 241396 370873
rect 241480 370813 241514 370873
rect 241638 370813 241672 370873
rect 241756 370813 241790 370873
rect 241914 370813 241948 370873
rect 242032 370813 242066 370873
rect 242190 370813 242224 370873
rect 242308 370813 242342 370873
rect 242466 370813 242500 370873
rect 242584 370813 242618 370873
rect 242742 370813 242776 370873
rect 242860 370813 242894 370873
rect 243018 370813 243052 370873
rect 243136 370813 243170 370873
rect 243294 370813 243328 370873
rect 243412 370813 243446 370873
rect 243570 370813 243604 370873
rect 243688 370813 243722 370873
rect 243846 370813 243880 370873
rect 243964 370813 243998 370873
rect 244122 370813 244156 370873
rect 244240 370813 244274 370873
rect 244398 370813 244432 370873
rect 244516 370813 244550 370873
rect 244674 370813 244708 370873
rect 244792 370813 244826 370873
rect 244950 370813 244984 370873
rect 245068 370813 245102 370873
rect 245226 370813 245260 370873
rect 245344 370813 245378 370873
rect 245502 370813 245536 370873
rect 245620 370813 245654 370873
rect 245778 370813 245812 370873
rect 245896 370813 245930 370873
rect 246054 370813 246088 370873
rect 246172 370813 246206 370873
rect 246330 370813 246364 370873
rect 246448 370813 246482 370873
rect 246606 370813 246640 370873
rect 58840 251371 58874 251431
rect 58998 251371 59032 251431
rect 59116 251371 59150 251431
rect 59274 251371 59308 251431
rect 59392 251371 59426 251431
rect 59550 251371 59584 251431
rect 59668 251371 59702 251431
rect 59826 251371 59860 251431
rect 59944 251371 59978 251431
rect 60102 251371 60136 251431
rect 147965 251495 147999 251555
rect 148123 251495 148157 251555
rect 148241 251495 148275 251555
rect 148399 251495 148433 251555
rect 148517 251495 148551 251555
rect 148675 251495 148709 251555
rect 148793 251495 148827 251555
rect 148951 251495 148985 251555
rect 149069 251495 149103 251555
rect 149227 251495 149261 251555
rect 149345 251495 149379 251555
rect 149503 251495 149537 251555
rect 149621 251495 149655 251555
rect 149779 251495 149813 251555
rect 149897 251495 149931 251555
rect 150055 251495 150089 251555
rect 150173 251495 150207 251555
rect 150331 251495 150365 251555
rect 150449 251495 150483 251555
rect 150607 251495 150641 251555
rect 234209 251695 234243 251755
rect 234367 251695 234401 251755
rect 234485 251695 234519 251755
rect 234643 251695 234677 251755
rect 234761 251695 234795 251755
rect 234919 251695 234953 251755
rect 235037 251695 235071 251755
rect 235195 251695 235229 251755
rect 235313 251695 235347 251755
rect 235471 251695 235505 251755
rect 235589 251695 235623 251755
rect 235747 251695 235781 251755
rect 235865 251695 235899 251755
rect 236023 251695 236057 251755
rect 236141 251695 236175 251755
rect 236299 251695 236333 251755
rect 236417 251695 236451 251755
rect 236575 251695 236609 251755
rect 236693 251695 236727 251755
rect 236851 251695 236885 251755
rect 236969 251695 237003 251755
rect 237127 251695 237161 251755
rect 237245 251695 237279 251755
rect 237403 251695 237437 251755
rect 237521 251695 237555 251755
rect 237679 251695 237713 251755
rect 237797 251695 237831 251755
rect 237955 251695 237989 251755
rect 238073 251695 238107 251755
rect 238231 251695 238265 251755
rect 238349 251695 238383 251755
rect 238507 251695 238541 251755
rect 238625 251695 238659 251755
rect 238783 251695 238817 251755
rect 238901 251695 238935 251755
rect 239059 251695 239093 251755
rect 239177 251695 239211 251755
rect 239335 251695 239369 251755
rect 239453 251695 239487 251755
rect 239611 251695 239645 251755
rect 239729 251695 239763 251755
rect 239887 251695 239921 251755
rect 240005 251695 240039 251755
rect 240163 251695 240197 251755
rect 240281 251695 240315 251755
rect 240439 251695 240473 251755
rect 240557 251695 240591 251755
rect 240715 251695 240749 251755
rect 240833 251695 240867 251755
rect 240991 251695 241025 251755
rect 241109 251695 241143 251755
rect 241267 251695 241301 251755
rect 241385 251695 241419 251755
rect 241543 251695 241577 251755
rect 241661 251695 241695 251755
rect 241819 251695 241853 251755
rect 241937 251695 241971 251755
rect 242095 251695 242129 251755
rect 242213 251695 242247 251755
rect 242371 251695 242405 251755
rect 242489 251695 242523 251755
rect 242647 251695 242681 251755
rect 242765 251695 242799 251755
rect 242923 251695 242957 251755
rect 243041 251695 243075 251755
rect 243199 251695 243233 251755
rect 243317 251695 243351 251755
rect 243475 251695 243509 251755
rect 243593 251695 243627 251755
rect 243751 251695 243785 251755
rect 243869 251695 243903 251755
rect 244027 251695 244061 251755
rect 244145 251695 244179 251755
rect 244303 251695 244337 251755
rect 244421 251695 244455 251755
rect 244579 251695 244613 251755
rect 244697 251695 244731 251755
rect 244855 251695 244889 251755
rect 244973 251695 245007 251755
rect 245131 251695 245165 251755
rect 245249 251695 245283 251755
rect 245407 251695 245441 251755
rect 245525 251695 245559 251755
rect 245683 251695 245717 251755
rect 245801 251695 245835 251755
rect 245959 251695 245993 251755
rect 246077 251695 246111 251755
rect 246235 251695 246269 251755
rect 246353 251695 246387 251755
rect 246511 251695 246545 251755
rect 246629 251695 246663 251755
rect 246787 251695 246821 251755
rect 246905 251695 246939 251755
rect 247063 251695 247097 251755
rect 247181 251695 247215 251755
rect 247339 251695 247373 251755
rect 247457 251695 247491 251755
rect 247615 251695 247649 251755
rect 247733 251695 247767 251755
rect 247891 251695 247925 251755
rect 248009 251695 248043 251755
rect 248167 251695 248201 251755
rect 413291 251409 413325 251469
rect 413449 251409 413483 251469
rect 413567 251409 413601 251469
rect 413725 251409 413759 251469
rect 413843 251409 413877 251469
rect 414001 251409 414035 251469
rect 414119 251409 414153 251469
rect 414277 251409 414311 251469
rect 414395 251409 414429 251469
rect 414553 251409 414587 251469
rect 414671 251409 414705 251469
rect 414829 251409 414863 251469
rect 414947 251409 414981 251469
rect 415105 251409 415139 251469
rect 415223 251409 415257 251469
rect 415381 251409 415415 251469
rect 415499 251409 415533 251469
rect 415657 251409 415691 251469
rect 415775 251409 415809 251469
rect 415933 251409 415967 251469
rect 416051 251409 416085 251469
rect 416209 251409 416243 251469
rect 416327 251409 416361 251469
rect 416485 251409 416519 251469
rect 416603 251409 416637 251469
rect 416761 251409 416795 251469
rect 416879 251409 416913 251469
rect 417037 251409 417071 251469
rect 417155 251409 417189 251469
rect 417313 251409 417347 251469
rect 417431 251409 417465 251469
rect 417589 251409 417623 251469
rect 417707 251409 417741 251469
rect 417865 251409 417899 251469
rect 417983 251409 418017 251469
rect 418141 251409 418175 251469
rect 418259 251409 418293 251469
rect 418417 251409 418451 251469
rect 418535 251409 418569 251469
rect 418693 251409 418727 251469
rect 418811 251409 418845 251469
rect 418969 251409 419003 251469
rect 419087 251409 419121 251469
rect 419245 251409 419279 251469
rect 419363 251409 419397 251469
rect 419521 251409 419555 251469
rect 419639 251409 419673 251469
rect 419797 251409 419831 251469
rect 419915 251409 419949 251469
rect 420073 251409 420107 251469
rect 420191 251409 420225 251469
rect 420349 251409 420383 251469
rect 420467 251409 420501 251469
rect 420625 251409 420659 251469
rect 420743 251409 420777 251469
rect 420901 251409 420935 251469
rect 421019 251409 421053 251469
rect 421177 251409 421211 251469
rect 421295 251409 421329 251469
rect 421453 251409 421487 251469
rect 421571 251409 421605 251469
rect 421729 251409 421763 251469
rect 421847 251409 421881 251469
rect 422005 251409 422039 251469
rect 422123 251409 422157 251469
rect 422281 251409 422315 251469
rect 422399 251409 422433 251469
rect 422557 251409 422591 251469
rect 422675 251409 422709 251469
rect 422833 251409 422867 251469
rect 422951 251409 422985 251469
rect 423109 251409 423143 251469
rect 423227 251409 423261 251469
rect 423385 251409 423419 251469
rect 423503 251409 423537 251469
rect 423661 251409 423695 251469
rect 423779 251409 423813 251469
rect 423937 251409 423971 251469
rect 424055 251409 424089 251469
rect 424213 251409 424247 251469
rect 424331 251409 424365 251469
rect 424489 251409 424523 251469
rect 424607 251409 424641 251469
rect 424765 251409 424799 251469
rect 424883 251409 424917 251469
rect 425041 251409 425075 251469
rect 425159 251409 425193 251469
rect 425317 251409 425351 251469
rect 425435 251409 425469 251469
rect 425593 251409 425627 251469
rect 425711 251409 425745 251469
rect 425869 251409 425903 251469
rect 425987 251409 426021 251469
rect 426145 251409 426179 251469
rect 426263 251409 426297 251469
rect 426421 251409 426455 251469
rect 426539 251409 426573 251469
rect 426697 251409 426731 251469
rect 426815 251409 426849 251469
rect 426973 251409 427007 251469
rect 427091 251409 427125 251469
rect 427249 251409 427283 251469
rect 503291 251409 503325 251469
rect 503449 251409 503483 251469
rect 503567 251409 503601 251469
rect 503725 251409 503759 251469
rect 503843 251409 503877 251469
rect 504001 251409 504035 251469
rect 504119 251409 504153 251469
rect 504277 251409 504311 251469
rect 504395 251409 504429 251469
rect 504553 251409 504587 251469
rect 504671 251409 504705 251469
rect 504829 251409 504863 251469
rect 504947 251409 504981 251469
rect 505105 251409 505139 251469
rect 505223 251409 505257 251469
rect 505381 251409 505415 251469
rect 505499 251409 505533 251469
rect 505657 251409 505691 251469
rect 505775 251409 505809 251469
rect 505933 251409 505967 251469
rect 506051 251409 506085 251469
rect 506209 251409 506243 251469
rect 506327 251409 506361 251469
rect 506485 251409 506519 251469
rect 506603 251409 506637 251469
rect 506761 251409 506795 251469
rect 506879 251409 506913 251469
rect 507037 251409 507071 251469
rect 507155 251409 507189 251469
rect 507313 251409 507347 251469
rect 507431 251409 507465 251469
rect 507589 251409 507623 251469
rect 507707 251409 507741 251469
rect 507865 251409 507899 251469
rect 507983 251409 508017 251469
rect 508141 251409 508175 251469
rect 508259 251409 508293 251469
rect 508417 251409 508451 251469
rect 508535 251409 508569 251469
rect 508693 251409 508727 251469
rect 508811 251409 508845 251469
rect 508969 251409 509003 251469
rect 509087 251409 509121 251469
rect 509245 251409 509279 251469
rect 509363 251409 509397 251469
rect 509521 251409 509555 251469
rect 509639 251409 509673 251469
rect 509797 251409 509831 251469
rect 509915 251409 509949 251469
rect 510073 251409 510107 251469
rect 510191 251409 510225 251469
rect 510349 251409 510383 251469
rect 510467 251409 510501 251469
rect 510625 251409 510659 251469
rect 510743 251409 510777 251469
rect 510901 251409 510935 251469
rect 511019 251409 511053 251469
rect 511177 251409 511211 251469
rect 511295 251409 511329 251469
rect 511453 251409 511487 251469
rect 511571 251409 511605 251469
rect 511729 251409 511763 251469
rect 511847 251409 511881 251469
rect 512005 251409 512039 251469
rect 512123 251409 512157 251469
rect 512281 251409 512315 251469
rect 512399 251409 512433 251469
rect 512557 251409 512591 251469
rect 512675 251409 512709 251469
rect 512833 251409 512867 251469
rect 512951 251409 512985 251469
rect 513109 251409 513143 251469
rect 513227 251409 513261 251469
rect 513385 251409 513419 251469
rect 513503 251409 513537 251469
rect 513661 251409 513695 251469
rect 513779 251409 513813 251469
rect 513937 251409 513971 251469
rect 514055 251409 514089 251469
rect 514213 251409 514247 251469
rect 514331 251409 514365 251469
rect 514489 251409 514523 251469
rect 514607 251409 514641 251469
rect 514765 251409 514799 251469
rect 514883 251409 514917 251469
rect 515041 251409 515075 251469
rect 515159 251409 515193 251469
rect 515317 251409 515351 251469
rect 515435 251409 515469 251469
rect 515593 251409 515627 251469
rect 515711 251409 515745 251469
rect 515869 251409 515903 251469
rect 515987 251409 516021 251469
rect 516145 251409 516179 251469
rect 516263 251409 516297 251469
rect 516421 251409 516455 251469
rect 516539 251409 516573 251469
rect 516697 251409 516731 251469
rect 516815 251409 516849 251469
rect 516973 251409 517007 251469
rect 517091 251409 517125 251469
rect 517249 251409 517283 251469
rect 322648 250813 322682 250873
rect 322806 250813 322840 250873
rect 322924 250813 322958 250873
rect 323082 250813 323116 250873
rect 323200 250813 323234 250873
rect 323358 250813 323392 250873
rect 323476 250813 323510 250873
rect 323634 250813 323668 250873
rect 323752 250813 323786 250873
rect 323910 250813 323944 250873
rect 324028 250813 324062 250873
rect 324186 250813 324220 250873
rect 324304 250813 324338 250873
rect 324462 250813 324496 250873
rect 324580 250813 324614 250873
rect 324738 250813 324772 250873
rect 324856 250813 324890 250873
rect 325014 250813 325048 250873
rect 325132 250813 325166 250873
rect 325290 250813 325324 250873
rect 325408 250813 325442 250873
rect 325566 250813 325600 250873
rect 325684 250813 325718 250873
rect 325842 250813 325876 250873
rect 325960 250813 325994 250873
rect 326118 250813 326152 250873
rect 326236 250813 326270 250873
rect 326394 250813 326428 250873
rect 326512 250813 326546 250873
rect 326670 250813 326704 250873
rect 326788 250813 326822 250873
rect 326946 250813 326980 250873
rect 327064 250813 327098 250873
rect 327222 250813 327256 250873
rect 327340 250813 327374 250873
rect 327498 250813 327532 250873
rect 327616 250813 327650 250873
rect 327774 250813 327808 250873
rect 327892 250813 327926 250873
rect 328050 250813 328084 250873
rect 328168 250813 328202 250873
rect 328326 250813 328360 250873
rect 328444 250813 328478 250873
rect 328602 250813 328636 250873
rect 328720 250813 328754 250873
rect 328878 250813 328912 250873
rect 328996 250813 329030 250873
rect 329154 250813 329188 250873
rect 329272 250813 329306 250873
rect 329430 250813 329464 250873
rect 329548 250813 329582 250873
rect 329706 250813 329740 250873
rect 329824 250813 329858 250873
rect 329982 250813 330016 250873
rect 330100 250813 330134 250873
rect 330258 250813 330292 250873
rect 330376 250813 330410 250873
rect 330534 250813 330568 250873
rect 330652 250813 330686 250873
rect 330810 250813 330844 250873
rect 330928 250813 330962 250873
rect 331086 250813 331120 250873
rect 331204 250813 331238 250873
rect 331362 250813 331396 250873
rect 331480 250813 331514 250873
rect 331638 250813 331672 250873
rect 331756 250813 331790 250873
rect 331914 250813 331948 250873
rect 332032 250813 332066 250873
rect 332190 250813 332224 250873
rect 332308 250813 332342 250873
rect 332466 250813 332500 250873
rect 332584 250813 332618 250873
rect 332742 250813 332776 250873
rect 332860 250813 332894 250873
rect 333018 250813 333052 250873
rect 333136 250813 333170 250873
rect 333294 250813 333328 250873
rect 333412 250813 333446 250873
rect 333570 250813 333604 250873
rect 333688 250813 333722 250873
rect 333846 250813 333880 250873
rect 333964 250813 333998 250873
rect 334122 250813 334156 250873
rect 334240 250813 334274 250873
rect 334398 250813 334432 250873
rect 334516 250813 334550 250873
rect 334674 250813 334708 250873
rect 334792 250813 334826 250873
rect 334950 250813 334984 250873
rect 335068 250813 335102 250873
rect 335226 250813 335260 250873
rect 335344 250813 335378 250873
rect 335502 250813 335536 250873
rect 335620 250813 335654 250873
rect 335778 250813 335812 250873
rect 335896 250813 335930 250873
rect 336054 250813 336088 250873
rect 336172 250813 336206 250873
rect 336330 250813 336364 250873
rect 336448 250813 336482 250873
rect 336606 250813 336640 250873
rect 149565 55795 149599 55971
rect 149723 55795 149757 55971
rect 239575 55505 239609 55681
rect 239733 55505 239767 55681
rect 419565 55795 419599 55971
rect 419723 55795 419757 55971
rect 509575 55505 509609 55681
rect 509733 55505 509767 55681
<< mvpdiffc >>
rect 419277 657278 419311 657454
rect 419435 657278 419469 657454
rect 329475 580354 329509 580530
rect 329633 580354 329667 580530
rect 149475 145354 149509 145530
rect 149633 145354 149667 145530
rect 419475 145354 419509 145530
rect 419633 145354 419667 145530
<< psubdiff >>
rect 329000 658048 329350 658082
rect 329000 657568 329034 658048
rect 329316 657986 329350 658048
rect 509000 658048 509350 658082
rect 329316 657568 329350 657630
rect 329000 657534 329350 657568
rect 509000 657568 509034 658048
rect 509316 657986 509350 658048
rect 509316 657568 509350 657630
rect 509000 657534 509350 657568
rect 149198 656124 149548 656158
rect 149198 655644 149232 656124
rect 149514 656062 149548 656124
rect 149514 655644 149548 655706
rect 149198 655610 149548 655644
rect 239198 581124 239548 581158
rect 239198 580644 239232 581124
rect 239514 581062 239548 581124
rect 239514 580644 239548 580706
rect 239198 580610 239548 580644
rect 239198 146124 239548 146158
rect 239198 145644 239232 146124
rect 239514 146062 239548 146124
rect 239514 145644 239548 145706
rect 239198 145610 239548 145644
rect 509198 146124 509548 146158
rect 509198 145644 509232 146124
rect 509514 146062 509548 146124
rect 509514 145644 509548 145706
rect 509198 145610 509548 145644
rect 59198 56124 59548 56158
rect 59198 55644 59232 56124
rect 59514 56062 59548 56124
rect 59514 55644 59548 55706
rect 59198 55610 59548 55644
rect 329198 56124 329548 56158
rect 329198 55644 329232 56124
rect 329514 56062 329548 56124
rect 329514 55644 329548 55706
rect 329198 55610 329548 55644
<< nsubdiff >>
rect 239181 656095 239531 656129
rect 239181 655597 239215 656095
rect 239497 656033 239531 656095
rect 239497 655597 239531 655659
rect 239181 655563 239531 655597
rect 59181 146095 59531 146129
rect 59181 145597 59215 146095
rect 59497 146033 59531 146095
rect 59497 145597 59531 145659
rect 59181 145563 59531 145597
rect 329181 146095 329531 146129
rect 329181 145597 329215 146095
rect 329497 146033 329531 146095
rect 329497 145597 329531 145659
rect 329181 145563 329531 145597
<< mvpsubdiff >>
rect 59419 656147 59903 656205
rect 59419 655619 59477 656147
rect 59845 656097 59903 656147
rect 59845 655669 59857 656097
rect 59891 655669 59903 656097
rect 59845 655619 59903 655669
rect 59419 655561 59903 655619
rect 419221 583071 419705 583129
rect 419221 582543 419279 583071
rect 419647 583021 419705 583071
rect 419647 582593 419659 583021
rect 419693 582593 419705 583021
rect 419647 582543 419705 582593
rect 419221 582485 419705 582543
rect 509231 582781 509715 582839
rect 509231 582253 509289 582781
rect 509657 582731 509715 582781
rect 509657 582303 509669 582731
rect 509703 582303 509715 582731
rect 509657 582253 509715 582303
rect 509231 582195 509715 582253
rect 59419 581147 59903 581205
rect 59419 580619 59477 581147
rect 59845 581097 59903 581147
rect 59845 580669 59857 581097
rect 59891 580669 59903 581097
rect 59845 580619 59903 580669
rect 59419 580561 59903 580619
rect 149429 580857 149913 580915
rect 149429 580329 149487 580857
rect 149855 580807 149913 580857
rect 149855 580379 149867 580807
rect 149901 580379 149913 580807
rect 149855 580329 149913 580379
rect 149429 580271 149913 580329
rect 323685 492323 337969 492381
rect 58695 491935 61663 491993
rect 58695 491523 58753 491935
rect 61605 491885 61663 491935
rect 61605 491573 61617 491885
rect 61651 491573 61663 491885
rect 323685 491911 323743 492323
rect 337911 492273 337969 492323
rect 337911 491961 337923 492273
rect 337957 491961 337969 492273
rect 337911 491911 337969 491961
rect 323685 491853 337969 491911
rect 508695 491935 511663 491993
rect 61605 491523 61663 491573
rect 58695 491465 61663 491523
rect 143145 491645 157429 491703
rect 143145 491233 143203 491645
rect 157371 491595 157429 491645
rect 157371 491283 157383 491595
rect 157417 491283 157429 491595
rect 157371 491233 157429 491283
rect 143145 491175 157429 491233
rect 418694 491607 420282 491665
rect 418694 491195 418752 491607
rect 420224 491557 420282 491607
rect 420224 491245 420236 491557
rect 420270 491245 420282 491557
rect 508695 491523 508753 491935
rect 511605 491885 511663 491935
rect 511605 491573 511617 491885
rect 511651 491573 511663 491885
rect 511605 491523 511663 491573
rect 508695 491465 511663 491523
rect 420224 491195 420282 491245
rect 418694 491137 420282 491195
rect 232502 491049 246786 491107
rect 232502 490637 232560 491049
rect 246728 490999 246786 491049
rect 246728 490687 246740 490999
rect 246774 490687 246786 490999
rect 246728 490637 246786 490687
rect 232502 490579 246786 490637
rect 323685 372323 337969 372381
rect 323685 371911 323743 372323
rect 337911 372273 337969 372323
rect 337911 371961 337923 372273
rect 337957 371961 337969 372273
rect 337911 371911 337969 371961
rect 323685 371853 337969 371911
rect 418695 371935 421663 371993
rect 53145 371645 67429 371703
rect 53145 371233 53203 371645
rect 67371 371595 67429 371645
rect 67371 371283 67383 371595
rect 67417 371283 67429 371595
rect 67371 371233 67429 371283
rect 53145 371175 67429 371233
rect 143145 371645 157429 371703
rect 143145 371233 143203 371645
rect 157371 371595 157429 371645
rect 157371 371283 157383 371595
rect 157417 371283 157429 371595
rect 418695 371523 418753 371935
rect 421605 371885 421663 371935
rect 421605 371573 421617 371885
rect 421651 371573 421663 371885
rect 421605 371523 421663 371573
rect 418695 371465 421663 371523
rect 508694 371607 510282 371665
rect 157371 371233 157429 371283
rect 143145 371175 157429 371233
rect 508694 371195 508752 371607
rect 510224 371557 510282 371607
rect 510224 371245 510236 371557
rect 510270 371245 510282 371557
rect 510224 371195 510282 371245
rect 508694 371137 510282 371195
rect 232502 371049 246786 371107
rect 232502 370637 232560 371049
rect 246728 370999 246786 371049
rect 246728 370687 246740 370999
rect 246774 370687 246786 370999
rect 246728 370637 246786 370687
rect 232502 370579 246786 370637
rect 234063 251931 248347 251989
rect 147819 251731 150787 251789
rect 58694 251607 60282 251665
rect 58694 251195 58752 251607
rect 60224 251557 60282 251607
rect 60224 251245 60236 251557
rect 60270 251245 60282 251557
rect 147819 251319 147877 251731
rect 150729 251681 150787 251731
rect 150729 251369 150741 251681
rect 150775 251369 150787 251681
rect 234063 251519 234121 251931
rect 248289 251881 248347 251931
rect 248289 251569 248301 251881
rect 248335 251569 248347 251881
rect 248289 251519 248347 251569
rect 234063 251461 248347 251519
rect 413145 251645 427429 251703
rect 150729 251319 150787 251369
rect 147819 251261 150787 251319
rect 60224 251195 60282 251245
rect 58694 251137 60282 251195
rect 413145 251233 413203 251645
rect 427371 251595 427429 251645
rect 427371 251283 427383 251595
rect 427417 251283 427429 251595
rect 427371 251233 427429 251283
rect 413145 251175 427429 251233
rect 503145 251645 517429 251703
rect 503145 251233 503203 251645
rect 517371 251595 517429 251645
rect 517371 251283 517383 251595
rect 517417 251283 517429 251595
rect 517371 251233 517429 251283
rect 503145 251175 517429 251233
rect 322502 251049 336786 251107
rect 322502 250637 322560 251049
rect 336728 250999 336786 251049
rect 336728 250687 336740 250999
rect 336774 250687 336786 250999
rect 336728 250637 336786 250687
rect 322502 250579 336786 250637
rect 149419 56147 149903 56205
rect 149419 55619 149477 56147
rect 149845 56097 149903 56147
rect 149845 55669 149857 56097
rect 149891 55669 149903 56097
rect 149845 55619 149903 55669
rect 149419 55561 149903 55619
rect 239429 55857 239913 55915
rect 239429 55329 239487 55857
rect 239855 55807 239913 55857
rect 239855 55379 239867 55807
rect 239901 55379 239913 55807
rect 419419 56147 419903 56205
rect 419419 55619 419477 56147
rect 419845 56097 419903 56147
rect 419845 55669 419857 56097
rect 419891 55669 419903 56097
rect 419845 55619 419903 55669
rect 419419 55561 419903 55619
rect 509429 55857 509913 55915
rect 239855 55329 239913 55379
rect 239429 55271 239913 55329
rect 509429 55329 509487 55857
rect 509855 55807 509913 55857
rect 509855 55379 509867 55807
rect 509901 55379 509913 55807
rect 509855 55329 509913 55379
rect 509429 55271 509913 55329
<< mvnsubdiff >>
rect 419131 657639 419615 657697
rect 419131 657093 419189 657639
rect 419557 657589 419615 657639
rect 419557 657143 419569 657589
rect 419603 657143 419615 657589
rect 419557 657093 419615 657143
rect 419131 657035 419615 657093
rect 329329 580715 329813 580773
rect 329329 580169 329387 580715
rect 329755 580665 329813 580715
rect 329755 580219 329767 580665
rect 329801 580219 329813 580665
rect 329755 580169 329813 580219
rect 329329 580111 329813 580169
rect 149329 145715 149813 145773
rect 149329 145169 149387 145715
rect 149755 145665 149813 145715
rect 149755 145219 149767 145665
rect 149801 145219 149813 145665
rect 419329 145715 419813 145773
rect 149755 145169 149813 145219
rect 149329 145111 149813 145169
rect 419329 145169 419387 145715
rect 419755 145665 419813 145715
rect 419755 145219 419767 145665
rect 419801 145219 419813 145665
rect 419755 145169 419813 145219
rect 419329 145111 419813 145169
<< psubdiffcont >>
rect 329316 657630 329350 657986
rect 509316 657630 509350 657986
rect 149514 655706 149548 656062
rect 239514 580706 239548 581062
rect 239514 145706 239548 146062
rect 509514 145706 509548 146062
rect 59514 55706 59548 56062
rect 329514 55706 329548 56062
<< nsubdiffcont >>
rect 239497 655659 239531 656033
rect 59497 145659 59531 146033
rect 329497 145659 329531 146033
<< mvpsubdiffcont >>
rect 59857 655669 59891 656097
rect 419659 582593 419693 583021
rect 509669 582303 509703 582731
rect 59857 580669 59891 581097
rect 149867 580379 149901 580807
rect 61617 491573 61651 491885
rect 337923 491961 337957 492273
rect 157383 491283 157417 491595
rect 420236 491245 420270 491557
rect 511617 491573 511651 491885
rect 246740 490687 246774 490999
rect 337923 371961 337957 372273
rect 67383 371283 67417 371595
rect 157383 371283 157417 371595
rect 421617 371573 421651 371885
rect 510236 371245 510270 371557
rect 246740 370687 246774 370999
rect 60236 251245 60270 251557
rect 150741 251369 150775 251681
rect 248301 251569 248335 251881
rect 427383 251283 427417 251595
rect 517383 251283 517417 251595
rect 336740 250687 336774 250999
rect 149857 55669 149891 56097
rect 239867 55379 239901 55807
rect 419857 55669 419891 56097
rect 509867 55379 509901 55807
<< mvnsubdiffcont >>
rect 419569 657143 419603 657589
rect 329767 580219 329801 580665
rect 149767 145219 149801 145665
rect 419767 145219 419801 145665
<< poly >>
rect 329142 657980 329208 657996
rect 329142 657946 329158 657980
rect 329192 657946 329208 657980
rect 329142 657930 329208 657946
rect 329160 657908 329190 657930
rect 329160 657686 329190 657708
rect 329142 657670 329208 657686
rect 329142 657636 329158 657670
rect 329192 657636 329208 657670
rect 329142 657620 329208 657636
rect 419323 657547 419423 657563
rect 419323 657513 419339 657547
rect 419407 657513 419423 657547
rect 419323 657466 419423 657513
rect 419323 657219 419423 657266
rect 419323 657185 419339 657219
rect 419407 657185 419423 657219
rect 419323 657169 419423 657185
rect 509142 657980 509208 657996
rect 509142 657946 509158 657980
rect 509192 657946 509208 657980
rect 509142 657930 509208 657946
rect 509160 657908 509190 657930
rect 509160 657686 509190 657708
rect 509142 657670 509208 657686
rect 509142 657636 509158 657670
rect 509192 657636 509208 657670
rect 509142 657620 509208 657636
rect 59611 656055 59711 656071
rect 59611 656021 59627 656055
rect 59695 656021 59711 656055
rect 59611 655983 59711 656021
rect 59611 655745 59711 655783
rect 59611 655711 59627 655745
rect 59695 655711 59711 655745
rect 59611 655695 59711 655711
rect 149340 656056 149406 656072
rect 149340 656022 149356 656056
rect 149390 656022 149406 656056
rect 149340 656006 149406 656022
rect 149358 655984 149388 656006
rect 149358 655762 149388 655784
rect 149340 655746 149406 655762
rect 149340 655712 149356 655746
rect 149390 655712 149406 655746
rect 149340 655696 149406 655712
rect 239323 656027 239389 656043
rect 239323 655993 239339 656027
rect 239373 655993 239389 656027
rect 239323 655977 239389 655993
rect 239341 655946 239371 655977
rect 239341 655715 239371 655746
rect 239323 655699 239389 655715
rect 239323 655665 239339 655699
rect 239373 655665 239389 655699
rect 239323 655649 239389 655665
rect 419413 582979 419513 582995
rect 419413 582945 419429 582979
rect 419497 582945 419513 582979
rect 419413 582907 419513 582945
rect 419413 582669 419513 582707
rect 419413 582635 419429 582669
rect 419497 582635 419513 582669
rect 419413 582619 419513 582635
rect 509423 582689 509523 582705
rect 509423 582655 509439 582689
rect 509507 582655 509523 582689
rect 509423 582617 509523 582655
rect 509423 582379 509523 582417
rect 509423 582345 509439 582379
rect 509507 582345 509523 582379
rect 509423 582329 509523 582345
rect 59611 581055 59711 581071
rect 59611 581021 59627 581055
rect 59695 581021 59711 581055
rect 59611 580983 59711 581021
rect 59611 580745 59711 580783
rect 59611 580711 59627 580745
rect 59695 580711 59711 580745
rect 59611 580695 59711 580711
rect 149621 580765 149721 580781
rect 149621 580731 149637 580765
rect 149705 580731 149721 580765
rect 149621 580693 149721 580731
rect 149621 580455 149721 580493
rect 149621 580421 149637 580455
rect 149705 580421 149721 580455
rect 149621 580405 149721 580421
rect 239340 581056 239406 581072
rect 239340 581022 239356 581056
rect 239390 581022 239406 581056
rect 239340 581006 239406 581022
rect 239358 580984 239388 581006
rect 239358 580762 239388 580784
rect 239340 580746 239406 580762
rect 239340 580712 239356 580746
rect 239390 580712 239406 580746
rect 239340 580696 239406 580712
rect 329521 580623 329621 580639
rect 329521 580589 329537 580623
rect 329605 580589 329621 580623
rect 329521 580542 329621 580589
rect 329521 580295 329621 580342
rect 329521 580261 329537 580295
rect 329605 580261 329621 580295
rect 329521 580245 329621 580261
rect 58887 491843 58987 491859
rect 58887 491809 58903 491843
rect 58971 491809 58987 491843
rect 58887 491771 58987 491809
rect 59163 491843 59263 491859
rect 59163 491809 59179 491843
rect 59247 491809 59263 491843
rect 59163 491771 59263 491809
rect 59439 491843 59539 491859
rect 59439 491809 59455 491843
rect 59523 491809 59539 491843
rect 59439 491771 59539 491809
rect 59715 491843 59815 491859
rect 59715 491809 59731 491843
rect 59799 491809 59815 491843
rect 59715 491771 59815 491809
rect 59991 491843 60091 491859
rect 59991 491809 60007 491843
rect 60075 491809 60091 491843
rect 59991 491771 60091 491809
rect 60267 491843 60367 491859
rect 60267 491809 60283 491843
rect 60351 491809 60367 491843
rect 60267 491771 60367 491809
rect 60543 491843 60643 491859
rect 60543 491809 60559 491843
rect 60627 491809 60643 491843
rect 60543 491771 60643 491809
rect 60819 491843 60919 491859
rect 60819 491809 60835 491843
rect 60903 491809 60919 491843
rect 60819 491771 60919 491809
rect 61095 491843 61195 491859
rect 61095 491809 61111 491843
rect 61179 491809 61195 491843
rect 61095 491771 61195 491809
rect 61371 491843 61471 491859
rect 61371 491809 61387 491843
rect 61455 491809 61471 491843
rect 61371 491771 61471 491809
rect 58887 491649 58987 491687
rect 58887 491615 58903 491649
rect 58971 491615 58987 491649
rect 58887 491599 58987 491615
rect 59163 491649 59263 491687
rect 59163 491615 59179 491649
rect 59247 491615 59263 491649
rect 59163 491599 59263 491615
rect 59439 491649 59539 491687
rect 59439 491615 59455 491649
rect 59523 491615 59539 491649
rect 59439 491599 59539 491615
rect 59715 491649 59815 491687
rect 59715 491615 59731 491649
rect 59799 491615 59815 491649
rect 59715 491599 59815 491615
rect 59991 491649 60091 491687
rect 59991 491615 60007 491649
rect 60075 491615 60091 491649
rect 59991 491599 60091 491615
rect 60267 491649 60367 491687
rect 60267 491615 60283 491649
rect 60351 491615 60367 491649
rect 60267 491599 60367 491615
rect 60543 491649 60643 491687
rect 60543 491615 60559 491649
rect 60627 491615 60643 491649
rect 60543 491599 60643 491615
rect 60819 491649 60919 491687
rect 60819 491615 60835 491649
rect 60903 491615 60919 491649
rect 60819 491599 60919 491615
rect 61095 491649 61195 491687
rect 61095 491615 61111 491649
rect 61179 491615 61195 491649
rect 61095 491599 61195 491615
rect 61371 491649 61471 491687
rect 61371 491615 61387 491649
rect 61455 491615 61471 491649
rect 61371 491599 61471 491615
rect 323877 492231 323977 492247
rect 323877 492197 323893 492231
rect 323961 492197 323977 492231
rect 323877 492159 323977 492197
rect 324153 492231 324253 492247
rect 324153 492197 324169 492231
rect 324237 492197 324253 492231
rect 324153 492159 324253 492197
rect 324429 492231 324529 492247
rect 324429 492197 324445 492231
rect 324513 492197 324529 492231
rect 324429 492159 324529 492197
rect 324705 492231 324805 492247
rect 324705 492197 324721 492231
rect 324789 492197 324805 492231
rect 324705 492159 324805 492197
rect 324981 492231 325081 492247
rect 324981 492197 324997 492231
rect 325065 492197 325081 492231
rect 324981 492159 325081 492197
rect 325257 492231 325357 492247
rect 325257 492197 325273 492231
rect 325341 492197 325357 492231
rect 325257 492159 325357 492197
rect 325533 492231 325633 492247
rect 325533 492197 325549 492231
rect 325617 492197 325633 492231
rect 325533 492159 325633 492197
rect 325809 492231 325909 492247
rect 325809 492197 325825 492231
rect 325893 492197 325909 492231
rect 325809 492159 325909 492197
rect 326085 492231 326185 492247
rect 326085 492197 326101 492231
rect 326169 492197 326185 492231
rect 326085 492159 326185 492197
rect 326361 492231 326461 492247
rect 326361 492197 326377 492231
rect 326445 492197 326461 492231
rect 326361 492159 326461 492197
rect 326637 492231 326737 492247
rect 326637 492197 326653 492231
rect 326721 492197 326737 492231
rect 326637 492159 326737 492197
rect 326913 492231 327013 492247
rect 326913 492197 326929 492231
rect 326997 492197 327013 492231
rect 326913 492159 327013 492197
rect 327189 492231 327289 492247
rect 327189 492197 327205 492231
rect 327273 492197 327289 492231
rect 327189 492159 327289 492197
rect 327465 492231 327565 492247
rect 327465 492197 327481 492231
rect 327549 492197 327565 492231
rect 327465 492159 327565 492197
rect 327741 492231 327841 492247
rect 327741 492197 327757 492231
rect 327825 492197 327841 492231
rect 327741 492159 327841 492197
rect 328017 492231 328117 492247
rect 328017 492197 328033 492231
rect 328101 492197 328117 492231
rect 328017 492159 328117 492197
rect 328293 492231 328393 492247
rect 328293 492197 328309 492231
rect 328377 492197 328393 492231
rect 328293 492159 328393 492197
rect 328569 492231 328669 492247
rect 328569 492197 328585 492231
rect 328653 492197 328669 492231
rect 328569 492159 328669 492197
rect 328845 492231 328945 492247
rect 328845 492197 328861 492231
rect 328929 492197 328945 492231
rect 328845 492159 328945 492197
rect 329121 492231 329221 492247
rect 329121 492197 329137 492231
rect 329205 492197 329221 492231
rect 329121 492159 329221 492197
rect 329397 492231 329497 492247
rect 329397 492197 329413 492231
rect 329481 492197 329497 492231
rect 329397 492159 329497 492197
rect 329673 492231 329773 492247
rect 329673 492197 329689 492231
rect 329757 492197 329773 492231
rect 329673 492159 329773 492197
rect 329949 492231 330049 492247
rect 329949 492197 329965 492231
rect 330033 492197 330049 492231
rect 329949 492159 330049 492197
rect 330225 492231 330325 492247
rect 330225 492197 330241 492231
rect 330309 492197 330325 492231
rect 330225 492159 330325 492197
rect 330501 492231 330601 492247
rect 330501 492197 330517 492231
rect 330585 492197 330601 492231
rect 330501 492159 330601 492197
rect 330777 492231 330877 492247
rect 330777 492197 330793 492231
rect 330861 492197 330877 492231
rect 330777 492159 330877 492197
rect 331053 492231 331153 492247
rect 331053 492197 331069 492231
rect 331137 492197 331153 492231
rect 331053 492159 331153 492197
rect 331329 492231 331429 492247
rect 331329 492197 331345 492231
rect 331413 492197 331429 492231
rect 331329 492159 331429 492197
rect 331605 492231 331705 492247
rect 331605 492197 331621 492231
rect 331689 492197 331705 492231
rect 331605 492159 331705 492197
rect 331881 492231 331981 492247
rect 331881 492197 331897 492231
rect 331965 492197 331981 492231
rect 331881 492159 331981 492197
rect 332157 492231 332257 492247
rect 332157 492197 332173 492231
rect 332241 492197 332257 492231
rect 332157 492159 332257 492197
rect 332433 492231 332533 492247
rect 332433 492197 332449 492231
rect 332517 492197 332533 492231
rect 332433 492159 332533 492197
rect 332709 492231 332809 492247
rect 332709 492197 332725 492231
rect 332793 492197 332809 492231
rect 332709 492159 332809 492197
rect 332985 492231 333085 492247
rect 332985 492197 333001 492231
rect 333069 492197 333085 492231
rect 332985 492159 333085 492197
rect 333261 492231 333361 492247
rect 333261 492197 333277 492231
rect 333345 492197 333361 492231
rect 333261 492159 333361 492197
rect 333537 492231 333637 492247
rect 333537 492197 333553 492231
rect 333621 492197 333637 492231
rect 333537 492159 333637 492197
rect 333813 492231 333913 492247
rect 333813 492197 333829 492231
rect 333897 492197 333913 492231
rect 333813 492159 333913 492197
rect 334089 492231 334189 492247
rect 334089 492197 334105 492231
rect 334173 492197 334189 492231
rect 334089 492159 334189 492197
rect 334365 492231 334465 492247
rect 334365 492197 334381 492231
rect 334449 492197 334465 492231
rect 334365 492159 334465 492197
rect 334641 492231 334741 492247
rect 334641 492197 334657 492231
rect 334725 492197 334741 492231
rect 334641 492159 334741 492197
rect 334917 492231 335017 492247
rect 334917 492197 334933 492231
rect 335001 492197 335017 492231
rect 334917 492159 335017 492197
rect 335193 492231 335293 492247
rect 335193 492197 335209 492231
rect 335277 492197 335293 492231
rect 335193 492159 335293 492197
rect 335469 492231 335569 492247
rect 335469 492197 335485 492231
rect 335553 492197 335569 492231
rect 335469 492159 335569 492197
rect 335745 492231 335845 492247
rect 335745 492197 335761 492231
rect 335829 492197 335845 492231
rect 335745 492159 335845 492197
rect 336021 492231 336121 492247
rect 336021 492197 336037 492231
rect 336105 492197 336121 492231
rect 336021 492159 336121 492197
rect 336297 492231 336397 492247
rect 336297 492197 336313 492231
rect 336381 492197 336397 492231
rect 336297 492159 336397 492197
rect 336573 492231 336673 492247
rect 336573 492197 336589 492231
rect 336657 492197 336673 492231
rect 336573 492159 336673 492197
rect 336849 492231 336949 492247
rect 336849 492197 336865 492231
rect 336933 492197 336949 492231
rect 336849 492159 336949 492197
rect 337125 492231 337225 492247
rect 337125 492197 337141 492231
rect 337209 492197 337225 492231
rect 337125 492159 337225 492197
rect 337401 492231 337501 492247
rect 337401 492197 337417 492231
rect 337485 492197 337501 492231
rect 337401 492159 337501 492197
rect 337677 492231 337777 492247
rect 337677 492197 337693 492231
rect 337761 492197 337777 492231
rect 337677 492159 337777 492197
rect 323877 492037 323977 492075
rect 323877 492003 323893 492037
rect 323961 492003 323977 492037
rect 323877 491987 323977 492003
rect 324153 492037 324253 492075
rect 324153 492003 324169 492037
rect 324237 492003 324253 492037
rect 324153 491987 324253 492003
rect 324429 492037 324529 492075
rect 324429 492003 324445 492037
rect 324513 492003 324529 492037
rect 324429 491987 324529 492003
rect 324705 492037 324805 492075
rect 324705 492003 324721 492037
rect 324789 492003 324805 492037
rect 324705 491987 324805 492003
rect 324981 492037 325081 492075
rect 324981 492003 324997 492037
rect 325065 492003 325081 492037
rect 324981 491987 325081 492003
rect 325257 492037 325357 492075
rect 325257 492003 325273 492037
rect 325341 492003 325357 492037
rect 325257 491987 325357 492003
rect 325533 492037 325633 492075
rect 325533 492003 325549 492037
rect 325617 492003 325633 492037
rect 325533 491987 325633 492003
rect 325809 492037 325909 492075
rect 325809 492003 325825 492037
rect 325893 492003 325909 492037
rect 325809 491987 325909 492003
rect 326085 492037 326185 492075
rect 326085 492003 326101 492037
rect 326169 492003 326185 492037
rect 326085 491987 326185 492003
rect 326361 492037 326461 492075
rect 326361 492003 326377 492037
rect 326445 492003 326461 492037
rect 326361 491987 326461 492003
rect 326637 492037 326737 492075
rect 326637 492003 326653 492037
rect 326721 492003 326737 492037
rect 326637 491987 326737 492003
rect 326913 492037 327013 492075
rect 326913 492003 326929 492037
rect 326997 492003 327013 492037
rect 326913 491987 327013 492003
rect 327189 492037 327289 492075
rect 327189 492003 327205 492037
rect 327273 492003 327289 492037
rect 327189 491987 327289 492003
rect 327465 492037 327565 492075
rect 327465 492003 327481 492037
rect 327549 492003 327565 492037
rect 327465 491987 327565 492003
rect 327741 492037 327841 492075
rect 327741 492003 327757 492037
rect 327825 492003 327841 492037
rect 327741 491987 327841 492003
rect 328017 492037 328117 492075
rect 328017 492003 328033 492037
rect 328101 492003 328117 492037
rect 328017 491987 328117 492003
rect 328293 492037 328393 492075
rect 328293 492003 328309 492037
rect 328377 492003 328393 492037
rect 328293 491987 328393 492003
rect 328569 492037 328669 492075
rect 328569 492003 328585 492037
rect 328653 492003 328669 492037
rect 328569 491987 328669 492003
rect 328845 492037 328945 492075
rect 328845 492003 328861 492037
rect 328929 492003 328945 492037
rect 328845 491987 328945 492003
rect 329121 492037 329221 492075
rect 329121 492003 329137 492037
rect 329205 492003 329221 492037
rect 329121 491987 329221 492003
rect 329397 492037 329497 492075
rect 329397 492003 329413 492037
rect 329481 492003 329497 492037
rect 329397 491987 329497 492003
rect 329673 492037 329773 492075
rect 329673 492003 329689 492037
rect 329757 492003 329773 492037
rect 329673 491987 329773 492003
rect 329949 492037 330049 492075
rect 329949 492003 329965 492037
rect 330033 492003 330049 492037
rect 329949 491987 330049 492003
rect 330225 492037 330325 492075
rect 330225 492003 330241 492037
rect 330309 492003 330325 492037
rect 330225 491987 330325 492003
rect 330501 492037 330601 492075
rect 330501 492003 330517 492037
rect 330585 492003 330601 492037
rect 330501 491987 330601 492003
rect 330777 492037 330877 492075
rect 330777 492003 330793 492037
rect 330861 492003 330877 492037
rect 330777 491987 330877 492003
rect 331053 492037 331153 492075
rect 331053 492003 331069 492037
rect 331137 492003 331153 492037
rect 331053 491987 331153 492003
rect 331329 492037 331429 492075
rect 331329 492003 331345 492037
rect 331413 492003 331429 492037
rect 331329 491987 331429 492003
rect 331605 492037 331705 492075
rect 331605 492003 331621 492037
rect 331689 492003 331705 492037
rect 331605 491987 331705 492003
rect 331881 492037 331981 492075
rect 331881 492003 331897 492037
rect 331965 492003 331981 492037
rect 331881 491987 331981 492003
rect 332157 492037 332257 492075
rect 332157 492003 332173 492037
rect 332241 492003 332257 492037
rect 332157 491987 332257 492003
rect 332433 492037 332533 492075
rect 332433 492003 332449 492037
rect 332517 492003 332533 492037
rect 332433 491987 332533 492003
rect 332709 492037 332809 492075
rect 332709 492003 332725 492037
rect 332793 492003 332809 492037
rect 332709 491987 332809 492003
rect 332985 492037 333085 492075
rect 332985 492003 333001 492037
rect 333069 492003 333085 492037
rect 332985 491987 333085 492003
rect 333261 492037 333361 492075
rect 333261 492003 333277 492037
rect 333345 492003 333361 492037
rect 333261 491987 333361 492003
rect 333537 492037 333637 492075
rect 333537 492003 333553 492037
rect 333621 492003 333637 492037
rect 333537 491987 333637 492003
rect 333813 492037 333913 492075
rect 333813 492003 333829 492037
rect 333897 492003 333913 492037
rect 333813 491987 333913 492003
rect 334089 492037 334189 492075
rect 334089 492003 334105 492037
rect 334173 492003 334189 492037
rect 334089 491987 334189 492003
rect 334365 492037 334465 492075
rect 334365 492003 334381 492037
rect 334449 492003 334465 492037
rect 334365 491987 334465 492003
rect 334641 492037 334741 492075
rect 334641 492003 334657 492037
rect 334725 492003 334741 492037
rect 334641 491987 334741 492003
rect 334917 492037 335017 492075
rect 334917 492003 334933 492037
rect 335001 492003 335017 492037
rect 334917 491987 335017 492003
rect 335193 492037 335293 492075
rect 335193 492003 335209 492037
rect 335277 492003 335293 492037
rect 335193 491987 335293 492003
rect 335469 492037 335569 492075
rect 335469 492003 335485 492037
rect 335553 492003 335569 492037
rect 335469 491987 335569 492003
rect 335745 492037 335845 492075
rect 335745 492003 335761 492037
rect 335829 492003 335845 492037
rect 335745 491987 335845 492003
rect 336021 492037 336121 492075
rect 336021 492003 336037 492037
rect 336105 492003 336121 492037
rect 336021 491987 336121 492003
rect 336297 492037 336397 492075
rect 336297 492003 336313 492037
rect 336381 492003 336397 492037
rect 336297 491987 336397 492003
rect 336573 492037 336673 492075
rect 336573 492003 336589 492037
rect 336657 492003 336673 492037
rect 336573 491987 336673 492003
rect 336849 492037 336949 492075
rect 336849 492003 336865 492037
rect 336933 492003 336949 492037
rect 336849 491987 336949 492003
rect 337125 492037 337225 492075
rect 337125 492003 337141 492037
rect 337209 492003 337225 492037
rect 337125 491987 337225 492003
rect 337401 492037 337501 492075
rect 337401 492003 337417 492037
rect 337485 492003 337501 492037
rect 337401 491987 337501 492003
rect 337677 492037 337777 492075
rect 337677 492003 337693 492037
rect 337761 492003 337777 492037
rect 337677 491987 337777 492003
rect 143337 491553 143437 491569
rect 143337 491519 143353 491553
rect 143421 491519 143437 491553
rect 143337 491481 143437 491519
rect 143613 491553 143713 491569
rect 143613 491519 143629 491553
rect 143697 491519 143713 491553
rect 143613 491481 143713 491519
rect 143889 491553 143989 491569
rect 143889 491519 143905 491553
rect 143973 491519 143989 491553
rect 143889 491481 143989 491519
rect 144165 491553 144265 491569
rect 144165 491519 144181 491553
rect 144249 491519 144265 491553
rect 144165 491481 144265 491519
rect 144441 491553 144541 491569
rect 144441 491519 144457 491553
rect 144525 491519 144541 491553
rect 144441 491481 144541 491519
rect 144717 491553 144817 491569
rect 144717 491519 144733 491553
rect 144801 491519 144817 491553
rect 144717 491481 144817 491519
rect 144993 491553 145093 491569
rect 144993 491519 145009 491553
rect 145077 491519 145093 491553
rect 144993 491481 145093 491519
rect 145269 491553 145369 491569
rect 145269 491519 145285 491553
rect 145353 491519 145369 491553
rect 145269 491481 145369 491519
rect 145545 491553 145645 491569
rect 145545 491519 145561 491553
rect 145629 491519 145645 491553
rect 145545 491481 145645 491519
rect 145821 491553 145921 491569
rect 145821 491519 145837 491553
rect 145905 491519 145921 491553
rect 145821 491481 145921 491519
rect 146097 491553 146197 491569
rect 146097 491519 146113 491553
rect 146181 491519 146197 491553
rect 146097 491481 146197 491519
rect 146373 491553 146473 491569
rect 146373 491519 146389 491553
rect 146457 491519 146473 491553
rect 146373 491481 146473 491519
rect 146649 491553 146749 491569
rect 146649 491519 146665 491553
rect 146733 491519 146749 491553
rect 146649 491481 146749 491519
rect 146925 491553 147025 491569
rect 146925 491519 146941 491553
rect 147009 491519 147025 491553
rect 146925 491481 147025 491519
rect 147201 491553 147301 491569
rect 147201 491519 147217 491553
rect 147285 491519 147301 491553
rect 147201 491481 147301 491519
rect 147477 491553 147577 491569
rect 147477 491519 147493 491553
rect 147561 491519 147577 491553
rect 147477 491481 147577 491519
rect 147753 491553 147853 491569
rect 147753 491519 147769 491553
rect 147837 491519 147853 491553
rect 147753 491481 147853 491519
rect 148029 491553 148129 491569
rect 148029 491519 148045 491553
rect 148113 491519 148129 491553
rect 148029 491481 148129 491519
rect 148305 491553 148405 491569
rect 148305 491519 148321 491553
rect 148389 491519 148405 491553
rect 148305 491481 148405 491519
rect 148581 491553 148681 491569
rect 148581 491519 148597 491553
rect 148665 491519 148681 491553
rect 148581 491481 148681 491519
rect 148857 491553 148957 491569
rect 148857 491519 148873 491553
rect 148941 491519 148957 491553
rect 148857 491481 148957 491519
rect 149133 491553 149233 491569
rect 149133 491519 149149 491553
rect 149217 491519 149233 491553
rect 149133 491481 149233 491519
rect 149409 491553 149509 491569
rect 149409 491519 149425 491553
rect 149493 491519 149509 491553
rect 149409 491481 149509 491519
rect 149685 491553 149785 491569
rect 149685 491519 149701 491553
rect 149769 491519 149785 491553
rect 149685 491481 149785 491519
rect 149961 491553 150061 491569
rect 149961 491519 149977 491553
rect 150045 491519 150061 491553
rect 149961 491481 150061 491519
rect 150237 491553 150337 491569
rect 150237 491519 150253 491553
rect 150321 491519 150337 491553
rect 150237 491481 150337 491519
rect 150513 491553 150613 491569
rect 150513 491519 150529 491553
rect 150597 491519 150613 491553
rect 150513 491481 150613 491519
rect 150789 491553 150889 491569
rect 150789 491519 150805 491553
rect 150873 491519 150889 491553
rect 150789 491481 150889 491519
rect 151065 491553 151165 491569
rect 151065 491519 151081 491553
rect 151149 491519 151165 491553
rect 151065 491481 151165 491519
rect 151341 491553 151441 491569
rect 151341 491519 151357 491553
rect 151425 491519 151441 491553
rect 151341 491481 151441 491519
rect 151617 491553 151717 491569
rect 151617 491519 151633 491553
rect 151701 491519 151717 491553
rect 151617 491481 151717 491519
rect 151893 491553 151993 491569
rect 151893 491519 151909 491553
rect 151977 491519 151993 491553
rect 151893 491481 151993 491519
rect 152169 491553 152269 491569
rect 152169 491519 152185 491553
rect 152253 491519 152269 491553
rect 152169 491481 152269 491519
rect 152445 491553 152545 491569
rect 152445 491519 152461 491553
rect 152529 491519 152545 491553
rect 152445 491481 152545 491519
rect 152721 491553 152821 491569
rect 152721 491519 152737 491553
rect 152805 491519 152821 491553
rect 152721 491481 152821 491519
rect 152997 491553 153097 491569
rect 152997 491519 153013 491553
rect 153081 491519 153097 491553
rect 152997 491481 153097 491519
rect 153273 491553 153373 491569
rect 153273 491519 153289 491553
rect 153357 491519 153373 491553
rect 153273 491481 153373 491519
rect 153549 491553 153649 491569
rect 153549 491519 153565 491553
rect 153633 491519 153649 491553
rect 153549 491481 153649 491519
rect 153825 491553 153925 491569
rect 153825 491519 153841 491553
rect 153909 491519 153925 491553
rect 153825 491481 153925 491519
rect 154101 491553 154201 491569
rect 154101 491519 154117 491553
rect 154185 491519 154201 491553
rect 154101 491481 154201 491519
rect 154377 491553 154477 491569
rect 154377 491519 154393 491553
rect 154461 491519 154477 491553
rect 154377 491481 154477 491519
rect 154653 491553 154753 491569
rect 154653 491519 154669 491553
rect 154737 491519 154753 491553
rect 154653 491481 154753 491519
rect 154929 491553 155029 491569
rect 154929 491519 154945 491553
rect 155013 491519 155029 491553
rect 154929 491481 155029 491519
rect 155205 491553 155305 491569
rect 155205 491519 155221 491553
rect 155289 491519 155305 491553
rect 155205 491481 155305 491519
rect 155481 491553 155581 491569
rect 155481 491519 155497 491553
rect 155565 491519 155581 491553
rect 155481 491481 155581 491519
rect 155757 491553 155857 491569
rect 155757 491519 155773 491553
rect 155841 491519 155857 491553
rect 155757 491481 155857 491519
rect 156033 491553 156133 491569
rect 156033 491519 156049 491553
rect 156117 491519 156133 491553
rect 156033 491481 156133 491519
rect 156309 491553 156409 491569
rect 156309 491519 156325 491553
rect 156393 491519 156409 491553
rect 156309 491481 156409 491519
rect 156585 491553 156685 491569
rect 156585 491519 156601 491553
rect 156669 491519 156685 491553
rect 156585 491481 156685 491519
rect 156861 491553 156961 491569
rect 156861 491519 156877 491553
rect 156945 491519 156961 491553
rect 156861 491481 156961 491519
rect 157137 491553 157237 491569
rect 157137 491519 157153 491553
rect 157221 491519 157237 491553
rect 157137 491481 157237 491519
rect 143337 491359 143437 491397
rect 143337 491325 143353 491359
rect 143421 491325 143437 491359
rect 143337 491309 143437 491325
rect 143613 491359 143713 491397
rect 143613 491325 143629 491359
rect 143697 491325 143713 491359
rect 143613 491309 143713 491325
rect 143889 491359 143989 491397
rect 143889 491325 143905 491359
rect 143973 491325 143989 491359
rect 143889 491309 143989 491325
rect 144165 491359 144265 491397
rect 144165 491325 144181 491359
rect 144249 491325 144265 491359
rect 144165 491309 144265 491325
rect 144441 491359 144541 491397
rect 144441 491325 144457 491359
rect 144525 491325 144541 491359
rect 144441 491309 144541 491325
rect 144717 491359 144817 491397
rect 144717 491325 144733 491359
rect 144801 491325 144817 491359
rect 144717 491309 144817 491325
rect 144993 491359 145093 491397
rect 144993 491325 145009 491359
rect 145077 491325 145093 491359
rect 144993 491309 145093 491325
rect 145269 491359 145369 491397
rect 145269 491325 145285 491359
rect 145353 491325 145369 491359
rect 145269 491309 145369 491325
rect 145545 491359 145645 491397
rect 145545 491325 145561 491359
rect 145629 491325 145645 491359
rect 145545 491309 145645 491325
rect 145821 491359 145921 491397
rect 145821 491325 145837 491359
rect 145905 491325 145921 491359
rect 145821 491309 145921 491325
rect 146097 491359 146197 491397
rect 146097 491325 146113 491359
rect 146181 491325 146197 491359
rect 146097 491309 146197 491325
rect 146373 491359 146473 491397
rect 146373 491325 146389 491359
rect 146457 491325 146473 491359
rect 146373 491309 146473 491325
rect 146649 491359 146749 491397
rect 146649 491325 146665 491359
rect 146733 491325 146749 491359
rect 146649 491309 146749 491325
rect 146925 491359 147025 491397
rect 146925 491325 146941 491359
rect 147009 491325 147025 491359
rect 146925 491309 147025 491325
rect 147201 491359 147301 491397
rect 147201 491325 147217 491359
rect 147285 491325 147301 491359
rect 147201 491309 147301 491325
rect 147477 491359 147577 491397
rect 147477 491325 147493 491359
rect 147561 491325 147577 491359
rect 147477 491309 147577 491325
rect 147753 491359 147853 491397
rect 147753 491325 147769 491359
rect 147837 491325 147853 491359
rect 147753 491309 147853 491325
rect 148029 491359 148129 491397
rect 148029 491325 148045 491359
rect 148113 491325 148129 491359
rect 148029 491309 148129 491325
rect 148305 491359 148405 491397
rect 148305 491325 148321 491359
rect 148389 491325 148405 491359
rect 148305 491309 148405 491325
rect 148581 491359 148681 491397
rect 148581 491325 148597 491359
rect 148665 491325 148681 491359
rect 148581 491309 148681 491325
rect 148857 491359 148957 491397
rect 148857 491325 148873 491359
rect 148941 491325 148957 491359
rect 148857 491309 148957 491325
rect 149133 491359 149233 491397
rect 149133 491325 149149 491359
rect 149217 491325 149233 491359
rect 149133 491309 149233 491325
rect 149409 491359 149509 491397
rect 149409 491325 149425 491359
rect 149493 491325 149509 491359
rect 149409 491309 149509 491325
rect 149685 491359 149785 491397
rect 149685 491325 149701 491359
rect 149769 491325 149785 491359
rect 149685 491309 149785 491325
rect 149961 491359 150061 491397
rect 149961 491325 149977 491359
rect 150045 491325 150061 491359
rect 149961 491309 150061 491325
rect 150237 491359 150337 491397
rect 150237 491325 150253 491359
rect 150321 491325 150337 491359
rect 150237 491309 150337 491325
rect 150513 491359 150613 491397
rect 150513 491325 150529 491359
rect 150597 491325 150613 491359
rect 150513 491309 150613 491325
rect 150789 491359 150889 491397
rect 150789 491325 150805 491359
rect 150873 491325 150889 491359
rect 150789 491309 150889 491325
rect 151065 491359 151165 491397
rect 151065 491325 151081 491359
rect 151149 491325 151165 491359
rect 151065 491309 151165 491325
rect 151341 491359 151441 491397
rect 151341 491325 151357 491359
rect 151425 491325 151441 491359
rect 151341 491309 151441 491325
rect 151617 491359 151717 491397
rect 151617 491325 151633 491359
rect 151701 491325 151717 491359
rect 151617 491309 151717 491325
rect 151893 491359 151993 491397
rect 151893 491325 151909 491359
rect 151977 491325 151993 491359
rect 151893 491309 151993 491325
rect 152169 491359 152269 491397
rect 152169 491325 152185 491359
rect 152253 491325 152269 491359
rect 152169 491309 152269 491325
rect 152445 491359 152545 491397
rect 152445 491325 152461 491359
rect 152529 491325 152545 491359
rect 152445 491309 152545 491325
rect 152721 491359 152821 491397
rect 152721 491325 152737 491359
rect 152805 491325 152821 491359
rect 152721 491309 152821 491325
rect 152997 491359 153097 491397
rect 152997 491325 153013 491359
rect 153081 491325 153097 491359
rect 152997 491309 153097 491325
rect 153273 491359 153373 491397
rect 153273 491325 153289 491359
rect 153357 491325 153373 491359
rect 153273 491309 153373 491325
rect 153549 491359 153649 491397
rect 153549 491325 153565 491359
rect 153633 491325 153649 491359
rect 153549 491309 153649 491325
rect 153825 491359 153925 491397
rect 153825 491325 153841 491359
rect 153909 491325 153925 491359
rect 153825 491309 153925 491325
rect 154101 491359 154201 491397
rect 154101 491325 154117 491359
rect 154185 491325 154201 491359
rect 154101 491309 154201 491325
rect 154377 491359 154477 491397
rect 154377 491325 154393 491359
rect 154461 491325 154477 491359
rect 154377 491309 154477 491325
rect 154653 491359 154753 491397
rect 154653 491325 154669 491359
rect 154737 491325 154753 491359
rect 154653 491309 154753 491325
rect 154929 491359 155029 491397
rect 154929 491325 154945 491359
rect 155013 491325 155029 491359
rect 154929 491309 155029 491325
rect 155205 491359 155305 491397
rect 155205 491325 155221 491359
rect 155289 491325 155305 491359
rect 155205 491309 155305 491325
rect 155481 491359 155581 491397
rect 155481 491325 155497 491359
rect 155565 491325 155581 491359
rect 155481 491309 155581 491325
rect 155757 491359 155857 491397
rect 155757 491325 155773 491359
rect 155841 491325 155857 491359
rect 155757 491309 155857 491325
rect 156033 491359 156133 491397
rect 156033 491325 156049 491359
rect 156117 491325 156133 491359
rect 156033 491309 156133 491325
rect 156309 491359 156409 491397
rect 156309 491325 156325 491359
rect 156393 491325 156409 491359
rect 156309 491309 156409 491325
rect 156585 491359 156685 491397
rect 156585 491325 156601 491359
rect 156669 491325 156685 491359
rect 156585 491309 156685 491325
rect 156861 491359 156961 491397
rect 156861 491325 156877 491359
rect 156945 491325 156961 491359
rect 156861 491309 156961 491325
rect 157137 491359 157237 491397
rect 157137 491325 157153 491359
rect 157221 491325 157237 491359
rect 157137 491309 157237 491325
rect 418886 491515 418986 491531
rect 418886 491481 418902 491515
rect 418970 491481 418986 491515
rect 418886 491443 418986 491481
rect 419162 491515 419262 491531
rect 419162 491481 419178 491515
rect 419246 491481 419262 491515
rect 419162 491443 419262 491481
rect 419438 491515 419538 491531
rect 419438 491481 419454 491515
rect 419522 491481 419538 491515
rect 419438 491443 419538 491481
rect 419714 491515 419814 491531
rect 419714 491481 419730 491515
rect 419798 491481 419814 491515
rect 419714 491443 419814 491481
rect 419990 491515 420090 491531
rect 419990 491481 420006 491515
rect 420074 491481 420090 491515
rect 419990 491443 420090 491481
rect 418886 491321 418986 491359
rect 418886 491287 418902 491321
rect 418970 491287 418986 491321
rect 418886 491271 418986 491287
rect 419162 491321 419262 491359
rect 419162 491287 419178 491321
rect 419246 491287 419262 491321
rect 419162 491271 419262 491287
rect 419438 491321 419538 491359
rect 419438 491287 419454 491321
rect 419522 491287 419538 491321
rect 419438 491271 419538 491287
rect 419714 491321 419814 491359
rect 419714 491287 419730 491321
rect 419798 491287 419814 491321
rect 419714 491271 419814 491287
rect 419990 491321 420090 491359
rect 419990 491287 420006 491321
rect 420074 491287 420090 491321
rect 419990 491271 420090 491287
rect 508887 491843 508987 491859
rect 508887 491809 508903 491843
rect 508971 491809 508987 491843
rect 508887 491771 508987 491809
rect 509163 491843 509263 491859
rect 509163 491809 509179 491843
rect 509247 491809 509263 491843
rect 509163 491771 509263 491809
rect 509439 491843 509539 491859
rect 509439 491809 509455 491843
rect 509523 491809 509539 491843
rect 509439 491771 509539 491809
rect 509715 491843 509815 491859
rect 509715 491809 509731 491843
rect 509799 491809 509815 491843
rect 509715 491771 509815 491809
rect 509991 491843 510091 491859
rect 509991 491809 510007 491843
rect 510075 491809 510091 491843
rect 509991 491771 510091 491809
rect 510267 491843 510367 491859
rect 510267 491809 510283 491843
rect 510351 491809 510367 491843
rect 510267 491771 510367 491809
rect 510543 491843 510643 491859
rect 510543 491809 510559 491843
rect 510627 491809 510643 491843
rect 510543 491771 510643 491809
rect 510819 491843 510919 491859
rect 510819 491809 510835 491843
rect 510903 491809 510919 491843
rect 510819 491771 510919 491809
rect 511095 491843 511195 491859
rect 511095 491809 511111 491843
rect 511179 491809 511195 491843
rect 511095 491771 511195 491809
rect 511371 491843 511471 491859
rect 511371 491809 511387 491843
rect 511455 491809 511471 491843
rect 511371 491771 511471 491809
rect 508887 491649 508987 491687
rect 508887 491615 508903 491649
rect 508971 491615 508987 491649
rect 508887 491599 508987 491615
rect 509163 491649 509263 491687
rect 509163 491615 509179 491649
rect 509247 491615 509263 491649
rect 509163 491599 509263 491615
rect 509439 491649 509539 491687
rect 509439 491615 509455 491649
rect 509523 491615 509539 491649
rect 509439 491599 509539 491615
rect 509715 491649 509815 491687
rect 509715 491615 509731 491649
rect 509799 491615 509815 491649
rect 509715 491599 509815 491615
rect 509991 491649 510091 491687
rect 509991 491615 510007 491649
rect 510075 491615 510091 491649
rect 509991 491599 510091 491615
rect 510267 491649 510367 491687
rect 510267 491615 510283 491649
rect 510351 491615 510367 491649
rect 510267 491599 510367 491615
rect 510543 491649 510643 491687
rect 510543 491615 510559 491649
rect 510627 491615 510643 491649
rect 510543 491599 510643 491615
rect 510819 491649 510919 491687
rect 510819 491615 510835 491649
rect 510903 491615 510919 491649
rect 510819 491599 510919 491615
rect 511095 491649 511195 491687
rect 511095 491615 511111 491649
rect 511179 491615 511195 491649
rect 511095 491599 511195 491615
rect 511371 491649 511471 491687
rect 511371 491615 511387 491649
rect 511455 491615 511471 491649
rect 511371 491599 511471 491615
rect 232694 490957 232794 490973
rect 232694 490923 232710 490957
rect 232778 490923 232794 490957
rect 232694 490885 232794 490923
rect 232970 490957 233070 490973
rect 232970 490923 232986 490957
rect 233054 490923 233070 490957
rect 232970 490885 233070 490923
rect 233246 490957 233346 490973
rect 233246 490923 233262 490957
rect 233330 490923 233346 490957
rect 233246 490885 233346 490923
rect 233522 490957 233622 490973
rect 233522 490923 233538 490957
rect 233606 490923 233622 490957
rect 233522 490885 233622 490923
rect 233798 490957 233898 490973
rect 233798 490923 233814 490957
rect 233882 490923 233898 490957
rect 233798 490885 233898 490923
rect 234074 490957 234174 490973
rect 234074 490923 234090 490957
rect 234158 490923 234174 490957
rect 234074 490885 234174 490923
rect 234350 490957 234450 490973
rect 234350 490923 234366 490957
rect 234434 490923 234450 490957
rect 234350 490885 234450 490923
rect 234626 490957 234726 490973
rect 234626 490923 234642 490957
rect 234710 490923 234726 490957
rect 234626 490885 234726 490923
rect 234902 490957 235002 490973
rect 234902 490923 234918 490957
rect 234986 490923 235002 490957
rect 234902 490885 235002 490923
rect 235178 490957 235278 490973
rect 235178 490923 235194 490957
rect 235262 490923 235278 490957
rect 235178 490885 235278 490923
rect 235454 490957 235554 490973
rect 235454 490923 235470 490957
rect 235538 490923 235554 490957
rect 235454 490885 235554 490923
rect 235730 490957 235830 490973
rect 235730 490923 235746 490957
rect 235814 490923 235830 490957
rect 235730 490885 235830 490923
rect 236006 490957 236106 490973
rect 236006 490923 236022 490957
rect 236090 490923 236106 490957
rect 236006 490885 236106 490923
rect 236282 490957 236382 490973
rect 236282 490923 236298 490957
rect 236366 490923 236382 490957
rect 236282 490885 236382 490923
rect 236558 490957 236658 490973
rect 236558 490923 236574 490957
rect 236642 490923 236658 490957
rect 236558 490885 236658 490923
rect 236834 490957 236934 490973
rect 236834 490923 236850 490957
rect 236918 490923 236934 490957
rect 236834 490885 236934 490923
rect 237110 490957 237210 490973
rect 237110 490923 237126 490957
rect 237194 490923 237210 490957
rect 237110 490885 237210 490923
rect 237386 490957 237486 490973
rect 237386 490923 237402 490957
rect 237470 490923 237486 490957
rect 237386 490885 237486 490923
rect 237662 490957 237762 490973
rect 237662 490923 237678 490957
rect 237746 490923 237762 490957
rect 237662 490885 237762 490923
rect 237938 490957 238038 490973
rect 237938 490923 237954 490957
rect 238022 490923 238038 490957
rect 237938 490885 238038 490923
rect 238214 490957 238314 490973
rect 238214 490923 238230 490957
rect 238298 490923 238314 490957
rect 238214 490885 238314 490923
rect 238490 490957 238590 490973
rect 238490 490923 238506 490957
rect 238574 490923 238590 490957
rect 238490 490885 238590 490923
rect 238766 490957 238866 490973
rect 238766 490923 238782 490957
rect 238850 490923 238866 490957
rect 238766 490885 238866 490923
rect 239042 490957 239142 490973
rect 239042 490923 239058 490957
rect 239126 490923 239142 490957
rect 239042 490885 239142 490923
rect 239318 490957 239418 490973
rect 239318 490923 239334 490957
rect 239402 490923 239418 490957
rect 239318 490885 239418 490923
rect 239594 490957 239694 490973
rect 239594 490923 239610 490957
rect 239678 490923 239694 490957
rect 239594 490885 239694 490923
rect 239870 490957 239970 490973
rect 239870 490923 239886 490957
rect 239954 490923 239970 490957
rect 239870 490885 239970 490923
rect 240146 490957 240246 490973
rect 240146 490923 240162 490957
rect 240230 490923 240246 490957
rect 240146 490885 240246 490923
rect 240422 490957 240522 490973
rect 240422 490923 240438 490957
rect 240506 490923 240522 490957
rect 240422 490885 240522 490923
rect 240698 490957 240798 490973
rect 240698 490923 240714 490957
rect 240782 490923 240798 490957
rect 240698 490885 240798 490923
rect 240974 490957 241074 490973
rect 240974 490923 240990 490957
rect 241058 490923 241074 490957
rect 240974 490885 241074 490923
rect 241250 490957 241350 490973
rect 241250 490923 241266 490957
rect 241334 490923 241350 490957
rect 241250 490885 241350 490923
rect 241526 490957 241626 490973
rect 241526 490923 241542 490957
rect 241610 490923 241626 490957
rect 241526 490885 241626 490923
rect 241802 490957 241902 490973
rect 241802 490923 241818 490957
rect 241886 490923 241902 490957
rect 241802 490885 241902 490923
rect 242078 490957 242178 490973
rect 242078 490923 242094 490957
rect 242162 490923 242178 490957
rect 242078 490885 242178 490923
rect 242354 490957 242454 490973
rect 242354 490923 242370 490957
rect 242438 490923 242454 490957
rect 242354 490885 242454 490923
rect 242630 490957 242730 490973
rect 242630 490923 242646 490957
rect 242714 490923 242730 490957
rect 242630 490885 242730 490923
rect 242906 490957 243006 490973
rect 242906 490923 242922 490957
rect 242990 490923 243006 490957
rect 242906 490885 243006 490923
rect 243182 490957 243282 490973
rect 243182 490923 243198 490957
rect 243266 490923 243282 490957
rect 243182 490885 243282 490923
rect 243458 490957 243558 490973
rect 243458 490923 243474 490957
rect 243542 490923 243558 490957
rect 243458 490885 243558 490923
rect 243734 490957 243834 490973
rect 243734 490923 243750 490957
rect 243818 490923 243834 490957
rect 243734 490885 243834 490923
rect 244010 490957 244110 490973
rect 244010 490923 244026 490957
rect 244094 490923 244110 490957
rect 244010 490885 244110 490923
rect 244286 490957 244386 490973
rect 244286 490923 244302 490957
rect 244370 490923 244386 490957
rect 244286 490885 244386 490923
rect 244562 490957 244662 490973
rect 244562 490923 244578 490957
rect 244646 490923 244662 490957
rect 244562 490885 244662 490923
rect 244838 490957 244938 490973
rect 244838 490923 244854 490957
rect 244922 490923 244938 490957
rect 244838 490885 244938 490923
rect 245114 490957 245214 490973
rect 245114 490923 245130 490957
rect 245198 490923 245214 490957
rect 245114 490885 245214 490923
rect 245390 490957 245490 490973
rect 245390 490923 245406 490957
rect 245474 490923 245490 490957
rect 245390 490885 245490 490923
rect 245666 490957 245766 490973
rect 245666 490923 245682 490957
rect 245750 490923 245766 490957
rect 245666 490885 245766 490923
rect 245942 490957 246042 490973
rect 245942 490923 245958 490957
rect 246026 490923 246042 490957
rect 245942 490885 246042 490923
rect 246218 490957 246318 490973
rect 246218 490923 246234 490957
rect 246302 490923 246318 490957
rect 246218 490885 246318 490923
rect 246494 490957 246594 490973
rect 246494 490923 246510 490957
rect 246578 490923 246594 490957
rect 246494 490885 246594 490923
rect 232694 490763 232794 490801
rect 232694 490729 232710 490763
rect 232778 490729 232794 490763
rect 232694 490713 232794 490729
rect 232970 490763 233070 490801
rect 232970 490729 232986 490763
rect 233054 490729 233070 490763
rect 232970 490713 233070 490729
rect 233246 490763 233346 490801
rect 233246 490729 233262 490763
rect 233330 490729 233346 490763
rect 233246 490713 233346 490729
rect 233522 490763 233622 490801
rect 233522 490729 233538 490763
rect 233606 490729 233622 490763
rect 233522 490713 233622 490729
rect 233798 490763 233898 490801
rect 233798 490729 233814 490763
rect 233882 490729 233898 490763
rect 233798 490713 233898 490729
rect 234074 490763 234174 490801
rect 234074 490729 234090 490763
rect 234158 490729 234174 490763
rect 234074 490713 234174 490729
rect 234350 490763 234450 490801
rect 234350 490729 234366 490763
rect 234434 490729 234450 490763
rect 234350 490713 234450 490729
rect 234626 490763 234726 490801
rect 234626 490729 234642 490763
rect 234710 490729 234726 490763
rect 234626 490713 234726 490729
rect 234902 490763 235002 490801
rect 234902 490729 234918 490763
rect 234986 490729 235002 490763
rect 234902 490713 235002 490729
rect 235178 490763 235278 490801
rect 235178 490729 235194 490763
rect 235262 490729 235278 490763
rect 235178 490713 235278 490729
rect 235454 490763 235554 490801
rect 235454 490729 235470 490763
rect 235538 490729 235554 490763
rect 235454 490713 235554 490729
rect 235730 490763 235830 490801
rect 235730 490729 235746 490763
rect 235814 490729 235830 490763
rect 235730 490713 235830 490729
rect 236006 490763 236106 490801
rect 236006 490729 236022 490763
rect 236090 490729 236106 490763
rect 236006 490713 236106 490729
rect 236282 490763 236382 490801
rect 236282 490729 236298 490763
rect 236366 490729 236382 490763
rect 236282 490713 236382 490729
rect 236558 490763 236658 490801
rect 236558 490729 236574 490763
rect 236642 490729 236658 490763
rect 236558 490713 236658 490729
rect 236834 490763 236934 490801
rect 236834 490729 236850 490763
rect 236918 490729 236934 490763
rect 236834 490713 236934 490729
rect 237110 490763 237210 490801
rect 237110 490729 237126 490763
rect 237194 490729 237210 490763
rect 237110 490713 237210 490729
rect 237386 490763 237486 490801
rect 237386 490729 237402 490763
rect 237470 490729 237486 490763
rect 237386 490713 237486 490729
rect 237662 490763 237762 490801
rect 237662 490729 237678 490763
rect 237746 490729 237762 490763
rect 237662 490713 237762 490729
rect 237938 490763 238038 490801
rect 237938 490729 237954 490763
rect 238022 490729 238038 490763
rect 237938 490713 238038 490729
rect 238214 490763 238314 490801
rect 238214 490729 238230 490763
rect 238298 490729 238314 490763
rect 238214 490713 238314 490729
rect 238490 490763 238590 490801
rect 238490 490729 238506 490763
rect 238574 490729 238590 490763
rect 238490 490713 238590 490729
rect 238766 490763 238866 490801
rect 238766 490729 238782 490763
rect 238850 490729 238866 490763
rect 238766 490713 238866 490729
rect 239042 490763 239142 490801
rect 239042 490729 239058 490763
rect 239126 490729 239142 490763
rect 239042 490713 239142 490729
rect 239318 490763 239418 490801
rect 239318 490729 239334 490763
rect 239402 490729 239418 490763
rect 239318 490713 239418 490729
rect 239594 490763 239694 490801
rect 239594 490729 239610 490763
rect 239678 490729 239694 490763
rect 239594 490713 239694 490729
rect 239870 490763 239970 490801
rect 239870 490729 239886 490763
rect 239954 490729 239970 490763
rect 239870 490713 239970 490729
rect 240146 490763 240246 490801
rect 240146 490729 240162 490763
rect 240230 490729 240246 490763
rect 240146 490713 240246 490729
rect 240422 490763 240522 490801
rect 240422 490729 240438 490763
rect 240506 490729 240522 490763
rect 240422 490713 240522 490729
rect 240698 490763 240798 490801
rect 240698 490729 240714 490763
rect 240782 490729 240798 490763
rect 240698 490713 240798 490729
rect 240974 490763 241074 490801
rect 240974 490729 240990 490763
rect 241058 490729 241074 490763
rect 240974 490713 241074 490729
rect 241250 490763 241350 490801
rect 241250 490729 241266 490763
rect 241334 490729 241350 490763
rect 241250 490713 241350 490729
rect 241526 490763 241626 490801
rect 241526 490729 241542 490763
rect 241610 490729 241626 490763
rect 241526 490713 241626 490729
rect 241802 490763 241902 490801
rect 241802 490729 241818 490763
rect 241886 490729 241902 490763
rect 241802 490713 241902 490729
rect 242078 490763 242178 490801
rect 242078 490729 242094 490763
rect 242162 490729 242178 490763
rect 242078 490713 242178 490729
rect 242354 490763 242454 490801
rect 242354 490729 242370 490763
rect 242438 490729 242454 490763
rect 242354 490713 242454 490729
rect 242630 490763 242730 490801
rect 242630 490729 242646 490763
rect 242714 490729 242730 490763
rect 242630 490713 242730 490729
rect 242906 490763 243006 490801
rect 242906 490729 242922 490763
rect 242990 490729 243006 490763
rect 242906 490713 243006 490729
rect 243182 490763 243282 490801
rect 243182 490729 243198 490763
rect 243266 490729 243282 490763
rect 243182 490713 243282 490729
rect 243458 490763 243558 490801
rect 243458 490729 243474 490763
rect 243542 490729 243558 490763
rect 243458 490713 243558 490729
rect 243734 490763 243834 490801
rect 243734 490729 243750 490763
rect 243818 490729 243834 490763
rect 243734 490713 243834 490729
rect 244010 490763 244110 490801
rect 244010 490729 244026 490763
rect 244094 490729 244110 490763
rect 244010 490713 244110 490729
rect 244286 490763 244386 490801
rect 244286 490729 244302 490763
rect 244370 490729 244386 490763
rect 244286 490713 244386 490729
rect 244562 490763 244662 490801
rect 244562 490729 244578 490763
rect 244646 490729 244662 490763
rect 244562 490713 244662 490729
rect 244838 490763 244938 490801
rect 244838 490729 244854 490763
rect 244922 490729 244938 490763
rect 244838 490713 244938 490729
rect 245114 490763 245214 490801
rect 245114 490729 245130 490763
rect 245198 490729 245214 490763
rect 245114 490713 245214 490729
rect 245390 490763 245490 490801
rect 245390 490729 245406 490763
rect 245474 490729 245490 490763
rect 245390 490713 245490 490729
rect 245666 490763 245766 490801
rect 245666 490729 245682 490763
rect 245750 490729 245766 490763
rect 245666 490713 245766 490729
rect 245942 490763 246042 490801
rect 245942 490729 245958 490763
rect 246026 490729 246042 490763
rect 245942 490713 246042 490729
rect 246218 490763 246318 490801
rect 246218 490729 246234 490763
rect 246302 490729 246318 490763
rect 246218 490713 246318 490729
rect 246494 490763 246594 490801
rect 246494 490729 246510 490763
rect 246578 490729 246594 490763
rect 246494 490713 246594 490729
rect 323877 372231 323977 372247
rect 323877 372197 323893 372231
rect 323961 372197 323977 372231
rect 323877 372159 323977 372197
rect 324153 372231 324253 372247
rect 324153 372197 324169 372231
rect 324237 372197 324253 372231
rect 324153 372159 324253 372197
rect 324429 372231 324529 372247
rect 324429 372197 324445 372231
rect 324513 372197 324529 372231
rect 324429 372159 324529 372197
rect 324705 372231 324805 372247
rect 324705 372197 324721 372231
rect 324789 372197 324805 372231
rect 324705 372159 324805 372197
rect 324981 372231 325081 372247
rect 324981 372197 324997 372231
rect 325065 372197 325081 372231
rect 324981 372159 325081 372197
rect 325257 372231 325357 372247
rect 325257 372197 325273 372231
rect 325341 372197 325357 372231
rect 325257 372159 325357 372197
rect 325533 372231 325633 372247
rect 325533 372197 325549 372231
rect 325617 372197 325633 372231
rect 325533 372159 325633 372197
rect 325809 372231 325909 372247
rect 325809 372197 325825 372231
rect 325893 372197 325909 372231
rect 325809 372159 325909 372197
rect 326085 372231 326185 372247
rect 326085 372197 326101 372231
rect 326169 372197 326185 372231
rect 326085 372159 326185 372197
rect 326361 372231 326461 372247
rect 326361 372197 326377 372231
rect 326445 372197 326461 372231
rect 326361 372159 326461 372197
rect 326637 372231 326737 372247
rect 326637 372197 326653 372231
rect 326721 372197 326737 372231
rect 326637 372159 326737 372197
rect 326913 372231 327013 372247
rect 326913 372197 326929 372231
rect 326997 372197 327013 372231
rect 326913 372159 327013 372197
rect 327189 372231 327289 372247
rect 327189 372197 327205 372231
rect 327273 372197 327289 372231
rect 327189 372159 327289 372197
rect 327465 372231 327565 372247
rect 327465 372197 327481 372231
rect 327549 372197 327565 372231
rect 327465 372159 327565 372197
rect 327741 372231 327841 372247
rect 327741 372197 327757 372231
rect 327825 372197 327841 372231
rect 327741 372159 327841 372197
rect 328017 372231 328117 372247
rect 328017 372197 328033 372231
rect 328101 372197 328117 372231
rect 328017 372159 328117 372197
rect 328293 372231 328393 372247
rect 328293 372197 328309 372231
rect 328377 372197 328393 372231
rect 328293 372159 328393 372197
rect 328569 372231 328669 372247
rect 328569 372197 328585 372231
rect 328653 372197 328669 372231
rect 328569 372159 328669 372197
rect 328845 372231 328945 372247
rect 328845 372197 328861 372231
rect 328929 372197 328945 372231
rect 328845 372159 328945 372197
rect 329121 372231 329221 372247
rect 329121 372197 329137 372231
rect 329205 372197 329221 372231
rect 329121 372159 329221 372197
rect 329397 372231 329497 372247
rect 329397 372197 329413 372231
rect 329481 372197 329497 372231
rect 329397 372159 329497 372197
rect 329673 372231 329773 372247
rect 329673 372197 329689 372231
rect 329757 372197 329773 372231
rect 329673 372159 329773 372197
rect 329949 372231 330049 372247
rect 329949 372197 329965 372231
rect 330033 372197 330049 372231
rect 329949 372159 330049 372197
rect 330225 372231 330325 372247
rect 330225 372197 330241 372231
rect 330309 372197 330325 372231
rect 330225 372159 330325 372197
rect 330501 372231 330601 372247
rect 330501 372197 330517 372231
rect 330585 372197 330601 372231
rect 330501 372159 330601 372197
rect 330777 372231 330877 372247
rect 330777 372197 330793 372231
rect 330861 372197 330877 372231
rect 330777 372159 330877 372197
rect 331053 372231 331153 372247
rect 331053 372197 331069 372231
rect 331137 372197 331153 372231
rect 331053 372159 331153 372197
rect 331329 372231 331429 372247
rect 331329 372197 331345 372231
rect 331413 372197 331429 372231
rect 331329 372159 331429 372197
rect 331605 372231 331705 372247
rect 331605 372197 331621 372231
rect 331689 372197 331705 372231
rect 331605 372159 331705 372197
rect 331881 372231 331981 372247
rect 331881 372197 331897 372231
rect 331965 372197 331981 372231
rect 331881 372159 331981 372197
rect 332157 372231 332257 372247
rect 332157 372197 332173 372231
rect 332241 372197 332257 372231
rect 332157 372159 332257 372197
rect 332433 372231 332533 372247
rect 332433 372197 332449 372231
rect 332517 372197 332533 372231
rect 332433 372159 332533 372197
rect 332709 372231 332809 372247
rect 332709 372197 332725 372231
rect 332793 372197 332809 372231
rect 332709 372159 332809 372197
rect 332985 372231 333085 372247
rect 332985 372197 333001 372231
rect 333069 372197 333085 372231
rect 332985 372159 333085 372197
rect 333261 372231 333361 372247
rect 333261 372197 333277 372231
rect 333345 372197 333361 372231
rect 333261 372159 333361 372197
rect 333537 372231 333637 372247
rect 333537 372197 333553 372231
rect 333621 372197 333637 372231
rect 333537 372159 333637 372197
rect 333813 372231 333913 372247
rect 333813 372197 333829 372231
rect 333897 372197 333913 372231
rect 333813 372159 333913 372197
rect 334089 372231 334189 372247
rect 334089 372197 334105 372231
rect 334173 372197 334189 372231
rect 334089 372159 334189 372197
rect 334365 372231 334465 372247
rect 334365 372197 334381 372231
rect 334449 372197 334465 372231
rect 334365 372159 334465 372197
rect 334641 372231 334741 372247
rect 334641 372197 334657 372231
rect 334725 372197 334741 372231
rect 334641 372159 334741 372197
rect 334917 372231 335017 372247
rect 334917 372197 334933 372231
rect 335001 372197 335017 372231
rect 334917 372159 335017 372197
rect 335193 372231 335293 372247
rect 335193 372197 335209 372231
rect 335277 372197 335293 372231
rect 335193 372159 335293 372197
rect 335469 372231 335569 372247
rect 335469 372197 335485 372231
rect 335553 372197 335569 372231
rect 335469 372159 335569 372197
rect 335745 372231 335845 372247
rect 335745 372197 335761 372231
rect 335829 372197 335845 372231
rect 335745 372159 335845 372197
rect 336021 372231 336121 372247
rect 336021 372197 336037 372231
rect 336105 372197 336121 372231
rect 336021 372159 336121 372197
rect 336297 372231 336397 372247
rect 336297 372197 336313 372231
rect 336381 372197 336397 372231
rect 336297 372159 336397 372197
rect 336573 372231 336673 372247
rect 336573 372197 336589 372231
rect 336657 372197 336673 372231
rect 336573 372159 336673 372197
rect 336849 372231 336949 372247
rect 336849 372197 336865 372231
rect 336933 372197 336949 372231
rect 336849 372159 336949 372197
rect 337125 372231 337225 372247
rect 337125 372197 337141 372231
rect 337209 372197 337225 372231
rect 337125 372159 337225 372197
rect 337401 372231 337501 372247
rect 337401 372197 337417 372231
rect 337485 372197 337501 372231
rect 337401 372159 337501 372197
rect 337677 372231 337777 372247
rect 337677 372197 337693 372231
rect 337761 372197 337777 372231
rect 337677 372159 337777 372197
rect 323877 372037 323977 372075
rect 323877 372003 323893 372037
rect 323961 372003 323977 372037
rect 323877 371987 323977 372003
rect 324153 372037 324253 372075
rect 324153 372003 324169 372037
rect 324237 372003 324253 372037
rect 324153 371987 324253 372003
rect 324429 372037 324529 372075
rect 324429 372003 324445 372037
rect 324513 372003 324529 372037
rect 324429 371987 324529 372003
rect 324705 372037 324805 372075
rect 324705 372003 324721 372037
rect 324789 372003 324805 372037
rect 324705 371987 324805 372003
rect 324981 372037 325081 372075
rect 324981 372003 324997 372037
rect 325065 372003 325081 372037
rect 324981 371987 325081 372003
rect 325257 372037 325357 372075
rect 325257 372003 325273 372037
rect 325341 372003 325357 372037
rect 325257 371987 325357 372003
rect 325533 372037 325633 372075
rect 325533 372003 325549 372037
rect 325617 372003 325633 372037
rect 325533 371987 325633 372003
rect 325809 372037 325909 372075
rect 325809 372003 325825 372037
rect 325893 372003 325909 372037
rect 325809 371987 325909 372003
rect 326085 372037 326185 372075
rect 326085 372003 326101 372037
rect 326169 372003 326185 372037
rect 326085 371987 326185 372003
rect 326361 372037 326461 372075
rect 326361 372003 326377 372037
rect 326445 372003 326461 372037
rect 326361 371987 326461 372003
rect 326637 372037 326737 372075
rect 326637 372003 326653 372037
rect 326721 372003 326737 372037
rect 326637 371987 326737 372003
rect 326913 372037 327013 372075
rect 326913 372003 326929 372037
rect 326997 372003 327013 372037
rect 326913 371987 327013 372003
rect 327189 372037 327289 372075
rect 327189 372003 327205 372037
rect 327273 372003 327289 372037
rect 327189 371987 327289 372003
rect 327465 372037 327565 372075
rect 327465 372003 327481 372037
rect 327549 372003 327565 372037
rect 327465 371987 327565 372003
rect 327741 372037 327841 372075
rect 327741 372003 327757 372037
rect 327825 372003 327841 372037
rect 327741 371987 327841 372003
rect 328017 372037 328117 372075
rect 328017 372003 328033 372037
rect 328101 372003 328117 372037
rect 328017 371987 328117 372003
rect 328293 372037 328393 372075
rect 328293 372003 328309 372037
rect 328377 372003 328393 372037
rect 328293 371987 328393 372003
rect 328569 372037 328669 372075
rect 328569 372003 328585 372037
rect 328653 372003 328669 372037
rect 328569 371987 328669 372003
rect 328845 372037 328945 372075
rect 328845 372003 328861 372037
rect 328929 372003 328945 372037
rect 328845 371987 328945 372003
rect 329121 372037 329221 372075
rect 329121 372003 329137 372037
rect 329205 372003 329221 372037
rect 329121 371987 329221 372003
rect 329397 372037 329497 372075
rect 329397 372003 329413 372037
rect 329481 372003 329497 372037
rect 329397 371987 329497 372003
rect 329673 372037 329773 372075
rect 329673 372003 329689 372037
rect 329757 372003 329773 372037
rect 329673 371987 329773 372003
rect 329949 372037 330049 372075
rect 329949 372003 329965 372037
rect 330033 372003 330049 372037
rect 329949 371987 330049 372003
rect 330225 372037 330325 372075
rect 330225 372003 330241 372037
rect 330309 372003 330325 372037
rect 330225 371987 330325 372003
rect 330501 372037 330601 372075
rect 330501 372003 330517 372037
rect 330585 372003 330601 372037
rect 330501 371987 330601 372003
rect 330777 372037 330877 372075
rect 330777 372003 330793 372037
rect 330861 372003 330877 372037
rect 330777 371987 330877 372003
rect 331053 372037 331153 372075
rect 331053 372003 331069 372037
rect 331137 372003 331153 372037
rect 331053 371987 331153 372003
rect 331329 372037 331429 372075
rect 331329 372003 331345 372037
rect 331413 372003 331429 372037
rect 331329 371987 331429 372003
rect 331605 372037 331705 372075
rect 331605 372003 331621 372037
rect 331689 372003 331705 372037
rect 331605 371987 331705 372003
rect 331881 372037 331981 372075
rect 331881 372003 331897 372037
rect 331965 372003 331981 372037
rect 331881 371987 331981 372003
rect 332157 372037 332257 372075
rect 332157 372003 332173 372037
rect 332241 372003 332257 372037
rect 332157 371987 332257 372003
rect 332433 372037 332533 372075
rect 332433 372003 332449 372037
rect 332517 372003 332533 372037
rect 332433 371987 332533 372003
rect 332709 372037 332809 372075
rect 332709 372003 332725 372037
rect 332793 372003 332809 372037
rect 332709 371987 332809 372003
rect 332985 372037 333085 372075
rect 332985 372003 333001 372037
rect 333069 372003 333085 372037
rect 332985 371987 333085 372003
rect 333261 372037 333361 372075
rect 333261 372003 333277 372037
rect 333345 372003 333361 372037
rect 333261 371987 333361 372003
rect 333537 372037 333637 372075
rect 333537 372003 333553 372037
rect 333621 372003 333637 372037
rect 333537 371987 333637 372003
rect 333813 372037 333913 372075
rect 333813 372003 333829 372037
rect 333897 372003 333913 372037
rect 333813 371987 333913 372003
rect 334089 372037 334189 372075
rect 334089 372003 334105 372037
rect 334173 372003 334189 372037
rect 334089 371987 334189 372003
rect 334365 372037 334465 372075
rect 334365 372003 334381 372037
rect 334449 372003 334465 372037
rect 334365 371987 334465 372003
rect 334641 372037 334741 372075
rect 334641 372003 334657 372037
rect 334725 372003 334741 372037
rect 334641 371987 334741 372003
rect 334917 372037 335017 372075
rect 334917 372003 334933 372037
rect 335001 372003 335017 372037
rect 334917 371987 335017 372003
rect 335193 372037 335293 372075
rect 335193 372003 335209 372037
rect 335277 372003 335293 372037
rect 335193 371987 335293 372003
rect 335469 372037 335569 372075
rect 335469 372003 335485 372037
rect 335553 372003 335569 372037
rect 335469 371987 335569 372003
rect 335745 372037 335845 372075
rect 335745 372003 335761 372037
rect 335829 372003 335845 372037
rect 335745 371987 335845 372003
rect 336021 372037 336121 372075
rect 336021 372003 336037 372037
rect 336105 372003 336121 372037
rect 336021 371987 336121 372003
rect 336297 372037 336397 372075
rect 336297 372003 336313 372037
rect 336381 372003 336397 372037
rect 336297 371987 336397 372003
rect 336573 372037 336673 372075
rect 336573 372003 336589 372037
rect 336657 372003 336673 372037
rect 336573 371987 336673 372003
rect 336849 372037 336949 372075
rect 336849 372003 336865 372037
rect 336933 372003 336949 372037
rect 336849 371987 336949 372003
rect 337125 372037 337225 372075
rect 337125 372003 337141 372037
rect 337209 372003 337225 372037
rect 337125 371987 337225 372003
rect 337401 372037 337501 372075
rect 337401 372003 337417 372037
rect 337485 372003 337501 372037
rect 337401 371987 337501 372003
rect 337677 372037 337777 372075
rect 337677 372003 337693 372037
rect 337761 372003 337777 372037
rect 337677 371987 337777 372003
rect 53337 371553 53437 371569
rect 53337 371519 53353 371553
rect 53421 371519 53437 371553
rect 53337 371481 53437 371519
rect 53613 371553 53713 371569
rect 53613 371519 53629 371553
rect 53697 371519 53713 371553
rect 53613 371481 53713 371519
rect 53889 371553 53989 371569
rect 53889 371519 53905 371553
rect 53973 371519 53989 371553
rect 53889 371481 53989 371519
rect 54165 371553 54265 371569
rect 54165 371519 54181 371553
rect 54249 371519 54265 371553
rect 54165 371481 54265 371519
rect 54441 371553 54541 371569
rect 54441 371519 54457 371553
rect 54525 371519 54541 371553
rect 54441 371481 54541 371519
rect 54717 371553 54817 371569
rect 54717 371519 54733 371553
rect 54801 371519 54817 371553
rect 54717 371481 54817 371519
rect 54993 371553 55093 371569
rect 54993 371519 55009 371553
rect 55077 371519 55093 371553
rect 54993 371481 55093 371519
rect 55269 371553 55369 371569
rect 55269 371519 55285 371553
rect 55353 371519 55369 371553
rect 55269 371481 55369 371519
rect 55545 371553 55645 371569
rect 55545 371519 55561 371553
rect 55629 371519 55645 371553
rect 55545 371481 55645 371519
rect 55821 371553 55921 371569
rect 55821 371519 55837 371553
rect 55905 371519 55921 371553
rect 55821 371481 55921 371519
rect 56097 371553 56197 371569
rect 56097 371519 56113 371553
rect 56181 371519 56197 371553
rect 56097 371481 56197 371519
rect 56373 371553 56473 371569
rect 56373 371519 56389 371553
rect 56457 371519 56473 371553
rect 56373 371481 56473 371519
rect 56649 371553 56749 371569
rect 56649 371519 56665 371553
rect 56733 371519 56749 371553
rect 56649 371481 56749 371519
rect 56925 371553 57025 371569
rect 56925 371519 56941 371553
rect 57009 371519 57025 371553
rect 56925 371481 57025 371519
rect 57201 371553 57301 371569
rect 57201 371519 57217 371553
rect 57285 371519 57301 371553
rect 57201 371481 57301 371519
rect 57477 371553 57577 371569
rect 57477 371519 57493 371553
rect 57561 371519 57577 371553
rect 57477 371481 57577 371519
rect 57753 371553 57853 371569
rect 57753 371519 57769 371553
rect 57837 371519 57853 371553
rect 57753 371481 57853 371519
rect 58029 371553 58129 371569
rect 58029 371519 58045 371553
rect 58113 371519 58129 371553
rect 58029 371481 58129 371519
rect 58305 371553 58405 371569
rect 58305 371519 58321 371553
rect 58389 371519 58405 371553
rect 58305 371481 58405 371519
rect 58581 371553 58681 371569
rect 58581 371519 58597 371553
rect 58665 371519 58681 371553
rect 58581 371481 58681 371519
rect 58857 371553 58957 371569
rect 58857 371519 58873 371553
rect 58941 371519 58957 371553
rect 58857 371481 58957 371519
rect 59133 371553 59233 371569
rect 59133 371519 59149 371553
rect 59217 371519 59233 371553
rect 59133 371481 59233 371519
rect 59409 371553 59509 371569
rect 59409 371519 59425 371553
rect 59493 371519 59509 371553
rect 59409 371481 59509 371519
rect 59685 371553 59785 371569
rect 59685 371519 59701 371553
rect 59769 371519 59785 371553
rect 59685 371481 59785 371519
rect 59961 371553 60061 371569
rect 59961 371519 59977 371553
rect 60045 371519 60061 371553
rect 59961 371481 60061 371519
rect 60237 371553 60337 371569
rect 60237 371519 60253 371553
rect 60321 371519 60337 371553
rect 60237 371481 60337 371519
rect 60513 371553 60613 371569
rect 60513 371519 60529 371553
rect 60597 371519 60613 371553
rect 60513 371481 60613 371519
rect 60789 371553 60889 371569
rect 60789 371519 60805 371553
rect 60873 371519 60889 371553
rect 60789 371481 60889 371519
rect 61065 371553 61165 371569
rect 61065 371519 61081 371553
rect 61149 371519 61165 371553
rect 61065 371481 61165 371519
rect 61341 371553 61441 371569
rect 61341 371519 61357 371553
rect 61425 371519 61441 371553
rect 61341 371481 61441 371519
rect 61617 371553 61717 371569
rect 61617 371519 61633 371553
rect 61701 371519 61717 371553
rect 61617 371481 61717 371519
rect 61893 371553 61993 371569
rect 61893 371519 61909 371553
rect 61977 371519 61993 371553
rect 61893 371481 61993 371519
rect 62169 371553 62269 371569
rect 62169 371519 62185 371553
rect 62253 371519 62269 371553
rect 62169 371481 62269 371519
rect 62445 371553 62545 371569
rect 62445 371519 62461 371553
rect 62529 371519 62545 371553
rect 62445 371481 62545 371519
rect 62721 371553 62821 371569
rect 62721 371519 62737 371553
rect 62805 371519 62821 371553
rect 62721 371481 62821 371519
rect 62997 371553 63097 371569
rect 62997 371519 63013 371553
rect 63081 371519 63097 371553
rect 62997 371481 63097 371519
rect 63273 371553 63373 371569
rect 63273 371519 63289 371553
rect 63357 371519 63373 371553
rect 63273 371481 63373 371519
rect 63549 371553 63649 371569
rect 63549 371519 63565 371553
rect 63633 371519 63649 371553
rect 63549 371481 63649 371519
rect 63825 371553 63925 371569
rect 63825 371519 63841 371553
rect 63909 371519 63925 371553
rect 63825 371481 63925 371519
rect 64101 371553 64201 371569
rect 64101 371519 64117 371553
rect 64185 371519 64201 371553
rect 64101 371481 64201 371519
rect 64377 371553 64477 371569
rect 64377 371519 64393 371553
rect 64461 371519 64477 371553
rect 64377 371481 64477 371519
rect 64653 371553 64753 371569
rect 64653 371519 64669 371553
rect 64737 371519 64753 371553
rect 64653 371481 64753 371519
rect 64929 371553 65029 371569
rect 64929 371519 64945 371553
rect 65013 371519 65029 371553
rect 64929 371481 65029 371519
rect 65205 371553 65305 371569
rect 65205 371519 65221 371553
rect 65289 371519 65305 371553
rect 65205 371481 65305 371519
rect 65481 371553 65581 371569
rect 65481 371519 65497 371553
rect 65565 371519 65581 371553
rect 65481 371481 65581 371519
rect 65757 371553 65857 371569
rect 65757 371519 65773 371553
rect 65841 371519 65857 371553
rect 65757 371481 65857 371519
rect 66033 371553 66133 371569
rect 66033 371519 66049 371553
rect 66117 371519 66133 371553
rect 66033 371481 66133 371519
rect 66309 371553 66409 371569
rect 66309 371519 66325 371553
rect 66393 371519 66409 371553
rect 66309 371481 66409 371519
rect 66585 371553 66685 371569
rect 66585 371519 66601 371553
rect 66669 371519 66685 371553
rect 66585 371481 66685 371519
rect 66861 371553 66961 371569
rect 66861 371519 66877 371553
rect 66945 371519 66961 371553
rect 66861 371481 66961 371519
rect 67137 371553 67237 371569
rect 67137 371519 67153 371553
rect 67221 371519 67237 371553
rect 67137 371481 67237 371519
rect 53337 371359 53437 371397
rect 53337 371325 53353 371359
rect 53421 371325 53437 371359
rect 53337 371309 53437 371325
rect 53613 371359 53713 371397
rect 53613 371325 53629 371359
rect 53697 371325 53713 371359
rect 53613 371309 53713 371325
rect 53889 371359 53989 371397
rect 53889 371325 53905 371359
rect 53973 371325 53989 371359
rect 53889 371309 53989 371325
rect 54165 371359 54265 371397
rect 54165 371325 54181 371359
rect 54249 371325 54265 371359
rect 54165 371309 54265 371325
rect 54441 371359 54541 371397
rect 54441 371325 54457 371359
rect 54525 371325 54541 371359
rect 54441 371309 54541 371325
rect 54717 371359 54817 371397
rect 54717 371325 54733 371359
rect 54801 371325 54817 371359
rect 54717 371309 54817 371325
rect 54993 371359 55093 371397
rect 54993 371325 55009 371359
rect 55077 371325 55093 371359
rect 54993 371309 55093 371325
rect 55269 371359 55369 371397
rect 55269 371325 55285 371359
rect 55353 371325 55369 371359
rect 55269 371309 55369 371325
rect 55545 371359 55645 371397
rect 55545 371325 55561 371359
rect 55629 371325 55645 371359
rect 55545 371309 55645 371325
rect 55821 371359 55921 371397
rect 55821 371325 55837 371359
rect 55905 371325 55921 371359
rect 55821 371309 55921 371325
rect 56097 371359 56197 371397
rect 56097 371325 56113 371359
rect 56181 371325 56197 371359
rect 56097 371309 56197 371325
rect 56373 371359 56473 371397
rect 56373 371325 56389 371359
rect 56457 371325 56473 371359
rect 56373 371309 56473 371325
rect 56649 371359 56749 371397
rect 56649 371325 56665 371359
rect 56733 371325 56749 371359
rect 56649 371309 56749 371325
rect 56925 371359 57025 371397
rect 56925 371325 56941 371359
rect 57009 371325 57025 371359
rect 56925 371309 57025 371325
rect 57201 371359 57301 371397
rect 57201 371325 57217 371359
rect 57285 371325 57301 371359
rect 57201 371309 57301 371325
rect 57477 371359 57577 371397
rect 57477 371325 57493 371359
rect 57561 371325 57577 371359
rect 57477 371309 57577 371325
rect 57753 371359 57853 371397
rect 57753 371325 57769 371359
rect 57837 371325 57853 371359
rect 57753 371309 57853 371325
rect 58029 371359 58129 371397
rect 58029 371325 58045 371359
rect 58113 371325 58129 371359
rect 58029 371309 58129 371325
rect 58305 371359 58405 371397
rect 58305 371325 58321 371359
rect 58389 371325 58405 371359
rect 58305 371309 58405 371325
rect 58581 371359 58681 371397
rect 58581 371325 58597 371359
rect 58665 371325 58681 371359
rect 58581 371309 58681 371325
rect 58857 371359 58957 371397
rect 58857 371325 58873 371359
rect 58941 371325 58957 371359
rect 58857 371309 58957 371325
rect 59133 371359 59233 371397
rect 59133 371325 59149 371359
rect 59217 371325 59233 371359
rect 59133 371309 59233 371325
rect 59409 371359 59509 371397
rect 59409 371325 59425 371359
rect 59493 371325 59509 371359
rect 59409 371309 59509 371325
rect 59685 371359 59785 371397
rect 59685 371325 59701 371359
rect 59769 371325 59785 371359
rect 59685 371309 59785 371325
rect 59961 371359 60061 371397
rect 59961 371325 59977 371359
rect 60045 371325 60061 371359
rect 59961 371309 60061 371325
rect 60237 371359 60337 371397
rect 60237 371325 60253 371359
rect 60321 371325 60337 371359
rect 60237 371309 60337 371325
rect 60513 371359 60613 371397
rect 60513 371325 60529 371359
rect 60597 371325 60613 371359
rect 60513 371309 60613 371325
rect 60789 371359 60889 371397
rect 60789 371325 60805 371359
rect 60873 371325 60889 371359
rect 60789 371309 60889 371325
rect 61065 371359 61165 371397
rect 61065 371325 61081 371359
rect 61149 371325 61165 371359
rect 61065 371309 61165 371325
rect 61341 371359 61441 371397
rect 61341 371325 61357 371359
rect 61425 371325 61441 371359
rect 61341 371309 61441 371325
rect 61617 371359 61717 371397
rect 61617 371325 61633 371359
rect 61701 371325 61717 371359
rect 61617 371309 61717 371325
rect 61893 371359 61993 371397
rect 61893 371325 61909 371359
rect 61977 371325 61993 371359
rect 61893 371309 61993 371325
rect 62169 371359 62269 371397
rect 62169 371325 62185 371359
rect 62253 371325 62269 371359
rect 62169 371309 62269 371325
rect 62445 371359 62545 371397
rect 62445 371325 62461 371359
rect 62529 371325 62545 371359
rect 62445 371309 62545 371325
rect 62721 371359 62821 371397
rect 62721 371325 62737 371359
rect 62805 371325 62821 371359
rect 62721 371309 62821 371325
rect 62997 371359 63097 371397
rect 62997 371325 63013 371359
rect 63081 371325 63097 371359
rect 62997 371309 63097 371325
rect 63273 371359 63373 371397
rect 63273 371325 63289 371359
rect 63357 371325 63373 371359
rect 63273 371309 63373 371325
rect 63549 371359 63649 371397
rect 63549 371325 63565 371359
rect 63633 371325 63649 371359
rect 63549 371309 63649 371325
rect 63825 371359 63925 371397
rect 63825 371325 63841 371359
rect 63909 371325 63925 371359
rect 63825 371309 63925 371325
rect 64101 371359 64201 371397
rect 64101 371325 64117 371359
rect 64185 371325 64201 371359
rect 64101 371309 64201 371325
rect 64377 371359 64477 371397
rect 64377 371325 64393 371359
rect 64461 371325 64477 371359
rect 64377 371309 64477 371325
rect 64653 371359 64753 371397
rect 64653 371325 64669 371359
rect 64737 371325 64753 371359
rect 64653 371309 64753 371325
rect 64929 371359 65029 371397
rect 64929 371325 64945 371359
rect 65013 371325 65029 371359
rect 64929 371309 65029 371325
rect 65205 371359 65305 371397
rect 65205 371325 65221 371359
rect 65289 371325 65305 371359
rect 65205 371309 65305 371325
rect 65481 371359 65581 371397
rect 65481 371325 65497 371359
rect 65565 371325 65581 371359
rect 65481 371309 65581 371325
rect 65757 371359 65857 371397
rect 65757 371325 65773 371359
rect 65841 371325 65857 371359
rect 65757 371309 65857 371325
rect 66033 371359 66133 371397
rect 66033 371325 66049 371359
rect 66117 371325 66133 371359
rect 66033 371309 66133 371325
rect 66309 371359 66409 371397
rect 66309 371325 66325 371359
rect 66393 371325 66409 371359
rect 66309 371309 66409 371325
rect 66585 371359 66685 371397
rect 66585 371325 66601 371359
rect 66669 371325 66685 371359
rect 66585 371309 66685 371325
rect 66861 371359 66961 371397
rect 66861 371325 66877 371359
rect 66945 371325 66961 371359
rect 66861 371309 66961 371325
rect 67137 371359 67237 371397
rect 67137 371325 67153 371359
rect 67221 371325 67237 371359
rect 67137 371309 67237 371325
rect 143337 371553 143437 371569
rect 143337 371519 143353 371553
rect 143421 371519 143437 371553
rect 143337 371481 143437 371519
rect 143613 371553 143713 371569
rect 143613 371519 143629 371553
rect 143697 371519 143713 371553
rect 143613 371481 143713 371519
rect 143889 371553 143989 371569
rect 143889 371519 143905 371553
rect 143973 371519 143989 371553
rect 143889 371481 143989 371519
rect 144165 371553 144265 371569
rect 144165 371519 144181 371553
rect 144249 371519 144265 371553
rect 144165 371481 144265 371519
rect 144441 371553 144541 371569
rect 144441 371519 144457 371553
rect 144525 371519 144541 371553
rect 144441 371481 144541 371519
rect 144717 371553 144817 371569
rect 144717 371519 144733 371553
rect 144801 371519 144817 371553
rect 144717 371481 144817 371519
rect 144993 371553 145093 371569
rect 144993 371519 145009 371553
rect 145077 371519 145093 371553
rect 144993 371481 145093 371519
rect 145269 371553 145369 371569
rect 145269 371519 145285 371553
rect 145353 371519 145369 371553
rect 145269 371481 145369 371519
rect 145545 371553 145645 371569
rect 145545 371519 145561 371553
rect 145629 371519 145645 371553
rect 145545 371481 145645 371519
rect 145821 371553 145921 371569
rect 145821 371519 145837 371553
rect 145905 371519 145921 371553
rect 145821 371481 145921 371519
rect 146097 371553 146197 371569
rect 146097 371519 146113 371553
rect 146181 371519 146197 371553
rect 146097 371481 146197 371519
rect 146373 371553 146473 371569
rect 146373 371519 146389 371553
rect 146457 371519 146473 371553
rect 146373 371481 146473 371519
rect 146649 371553 146749 371569
rect 146649 371519 146665 371553
rect 146733 371519 146749 371553
rect 146649 371481 146749 371519
rect 146925 371553 147025 371569
rect 146925 371519 146941 371553
rect 147009 371519 147025 371553
rect 146925 371481 147025 371519
rect 147201 371553 147301 371569
rect 147201 371519 147217 371553
rect 147285 371519 147301 371553
rect 147201 371481 147301 371519
rect 147477 371553 147577 371569
rect 147477 371519 147493 371553
rect 147561 371519 147577 371553
rect 147477 371481 147577 371519
rect 147753 371553 147853 371569
rect 147753 371519 147769 371553
rect 147837 371519 147853 371553
rect 147753 371481 147853 371519
rect 148029 371553 148129 371569
rect 148029 371519 148045 371553
rect 148113 371519 148129 371553
rect 148029 371481 148129 371519
rect 148305 371553 148405 371569
rect 148305 371519 148321 371553
rect 148389 371519 148405 371553
rect 148305 371481 148405 371519
rect 148581 371553 148681 371569
rect 148581 371519 148597 371553
rect 148665 371519 148681 371553
rect 148581 371481 148681 371519
rect 148857 371553 148957 371569
rect 148857 371519 148873 371553
rect 148941 371519 148957 371553
rect 148857 371481 148957 371519
rect 149133 371553 149233 371569
rect 149133 371519 149149 371553
rect 149217 371519 149233 371553
rect 149133 371481 149233 371519
rect 149409 371553 149509 371569
rect 149409 371519 149425 371553
rect 149493 371519 149509 371553
rect 149409 371481 149509 371519
rect 149685 371553 149785 371569
rect 149685 371519 149701 371553
rect 149769 371519 149785 371553
rect 149685 371481 149785 371519
rect 149961 371553 150061 371569
rect 149961 371519 149977 371553
rect 150045 371519 150061 371553
rect 149961 371481 150061 371519
rect 150237 371553 150337 371569
rect 150237 371519 150253 371553
rect 150321 371519 150337 371553
rect 150237 371481 150337 371519
rect 150513 371553 150613 371569
rect 150513 371519 150529 371553
rect 150597 371519 150613 371553
rect 150513 371481 150613 371519
rect 150789 371553 150889 371569
rect 150789 371519 150805 371553
rect 150873 371519 150889 371553
rect 150789 371481 150889 371519
rect 151065 371553 151165 371569
rect 151065 371519 151081 371553
rect 151149 371519 151165 371553
rect 151065 371481 151165 371519
rect 151341 371553 151441 371569
rect 151341 371519 151357 371553
rect 151425 371519 151441 371553
rect 151341 371481 151441 371519
rect 151617 371553 151717 371569
rect 151617 371519 151633 371553
rect 151701 371519 151717 371553
rect 151617 371481 151717 371519
rect 151893 371553 151993 371569
rect 151893 371519 151909 371553
rect 151977 371519 151993 371553
rect 151893 371481 151993 371519
rect 152169 371553 152269 371569
rect 152169 371519 152185 371553
rect 152253 371519 152269 371553
rect 152169 371481 152269 371519
rect 152445 371553 152545 371569
rect 152445 371519 152461 371553
rect 152529 371519 152545 371553
rect 152445 371481 152545 371519
rect 152721 371553 152821 371569
rect 152721 371519 152737 371553
rect 152805 371519 152821 371553
rect 152721 371481 152821 371519
rect 152997 371553 153097 371569
rect 152997 371519 153013 371553
rect 153081 371519 153097 371553
rect 152997 371481 153097 371519
rect 153273 371553 153373 371569
rect 153273 371519 153289 371553
rect 153357 371519 153373 371553
rect 153273 371481 153373 371519
rect 153549 371553 153649 371569
rect 153549 371519 153565 371553
rect 153633 371519 153649 371553
rect 153549 371481 153649 371519
rect 153825 371553 153925 371569
rect 153825 371519 153841 371553
rect 153909 371519 153925 371553
rect 153825 371481 153925 371519
rect 154101 371553 154201 371569
rect 154101 371519 154117 371553
rect 154185 371519 154201 371553
rect 154101 371481 154201 371519
rect 154377 371553 154477 371569
rect 154377 371519 154393 371553
rect 154461 371519 154477 371553
rect 154377 371481 154477 371519
rect 154653 371553 154753 371569
rect 154653 371519 154669 371553
rect 154737 371519 154753 371553
rect 154653 371481 154753 371519
rect 154929 371553 155029 371569
rect 154929 371519 154945 371553
rect 155013 371519 155029 371553
rect 154929 371481 155029 371519
rect 155205 371553 155305 371569
rect 155205 371519 155221 371553
rect 155289 371519 155305 371553
rect 155205 371481 155305 371519
rect 155481 371553 155581 371569
rect 155481 371519 155497 371553
rect 155565 371519 155581 371553
rect 155481 371481 155581 371519
rect 155757 371553 155857 371569
rect 155757 371519 155773 371553
rect 155841 371519 155857 371553
rect 155757 371481 155857 371519
rect 156033 371553 156133 371569
rect 156033 371519 156049 371553
rect 156117 371519 156133 371553
rect 156033 371481 156133 371519
rect 156309 371553 156409 371569
rect 156309 371519 156325 371553
rect 156393 371519 156409 371553
rect 156309 371481 156409 371519
rect 156585 371553 156685 371569
rect 156585 371519 156601 371553
rect 156669 371519 156685 371553
rect 156585 371481 156685 371519
rect 156861 371553 156961 371569
rect 156861 371519 156877 371553
rect 156945 371519 156961 371553
rect 156861 371481 156961 371519
rect 157137 371553 157237 371569
rect 157137 371519 157153 371553
rect 157221 371519 157237 371553
rect 157137 371481 157237 371519
rect 143337 371359 143437 371397
rect 143337 371325 143353 371359
rect 143421 371325 143437 371359
rect 143337 371309 143437 371325
rect 143613 371359 143713 371397
rect 143613 371325 143629 371359
rect 143697 371325 143713 371359
rect 143613 371309 143713 371325
rect 143889 371359 143989 371397
rect 143889 371325 143905 371359
rect 143973 371325 143989 371359
rect 143889 371309 143989 371325
rect 144165 371359 144265 371397
rect 144165 371325 144181 371359
rect 144249 371325 144265 371359
rect 144165 371309 144265 371325
rect 144441 371359 144541 371397
rect 144441 371325 144457 371359
rect 144525 371325 144541 371359
rect 144441 371309 144541 371325
rect 144717 371359 144817 371397
rect 144717 371325 144733 371359
rect 144801 371325 144817 371359
rect 144717 371309 144817 371325
rect 144993 371359 145093 371397
rect 144993 371325 145009 371359
rect 145077 371325 145093 371359
rect 144993 371309 145093 371325
rect 145269 371359 145369 371397
rect 145269 371325 145285 371359
rect 145353 371325 145369 371359
rect 145269 371309 145369 371325
rect 145545 371359 145645 371397
rect 145545 371325 145561 371359
rect 145629 371325 145645 371359
rect 145545 371309 145645 371325
rect 145821 371359 145921 371397
rect 145821 371325 145837 371359
rect 145905 371325 145921 371359
rect 145821 371309 145921 371325
rect 146097 371359 146197 371397
rect 146097 371325 146113 371359
rect 146181 371325 146197 371359
rect 146097 371309 146197 371325
rect 146373 371359 146473 371397
rect 146373 371325 146389 371359
rect 146457 371325 146473 371359
rect 146373 371309 146473 371325
rect 146649 371359 146749 371397
rect 146649 371325 146665 371359
rect 146733 371325 146749 371359
rect 146649 371309 146749 371325
rect 146925 371359 147025 371397
rect 146925 371325 146941 371359
rect 147009 371325 147025 371359
rect 146925 371309 147025 371325
rect 147201 371359 147301 371397
rect 147201 371325 147217 371359
rect 147285 371325 147301 371359
rect 147201 371309 147301 371325
rect 147477 371359 147577 371397
rect 147477 371325 147493 371359
rect 147561 371325 147577 371359
rect 147477 371309 147577 371325
rect 147753 371359 147853 371397
rect 147753 371325 147769 371359
rect 147837 371325 147853 371359
rect 147753 371309 147853 371325
rect 148029 371359 148129 371397
rect 148029 371325 148045 371359
rect 148113 371325 148129 371359
rect 148029 371309 148129 371325
rect 148305 371359 148405 371397
rect 148305 371325 148321 371359
rect 148389 371325 148405 371359
rect 148305 371309 148405 371325
rect 148581 371359 148681 371397
rect 148581 371325 148597 371359
rect 148665 371325 148681 371359
rect 148581 371309 148681 371325
rect 148857 371359 148957 371397
rect 148857 371325 148873 371359
rect 148941 371325 148957 371359
rect 148857 371309 148957 371325
rect 149133 371359 149233 371397
rect 149133 371325 149149 371359
rect 149217 371325 149233 371359
rect 149133 371309 149233 371325
rect 149409 371359 149509 371397
rect 149409 371325 149425 371359
rect 149493 371325 149509 371359
rect 149409 371309 149509 371325
rect 149685 371359 149785 371397
rect 149685 371325 149701 371359
rect 149769 371325 149785 371359
rect 149685 371309 149785 371325
rect 149961 371359 150061 371397
rect 149961 371325 149977 371359
rect 150045 371325 150061 371359
rect 149961 371309 150061 371325
rect 150237 371359 150337 371397
rect 150237 371325 150253 371359
rect 150321 371325 150337 371359
rect 150237 371309 150337 371325
rect 150513 371359 150613 371397
rect 150513 371325 150529 371359
rect 150597 371325 150613 371359
rect 150513 371309 150613 371325
rect 150789 371359 150889 371397
rect 150789 371325 150805 371359
rect 150873 371325 150889 371359
rect 150789 371309 150889 371325
rect 151065 371359 151165 371397
rect 151065 371325 151081 371359
rect 151149 371325 151165 371359
rect 151065 371309 151165 371325
rect 151341 371359 151441 371397
rect 151341 371325 151357 371359
rect 151425 371325 151441 371359
rect 151341 371309 151441 371325
rect 151617 371359 151717 371397
rect 151617 371325 151633 371359
rect 151701 371325 151717 371359
rect 151617 371309 151717 371325
rect 151893 371359 151993 371397
rect 151893 371325 151909 371359
rect 151977 371325 151993 371359
rect 151893 371309 151993 371325
rect 152169 371359 152269 371397
rect 152169 371325 152185 371359
rect 152253 371325 152269 371359
rect 152169 371309 152269 371325
rect 152445 371359 152545 371397
rect 152445 371325 152461 371359
rect 152529 371325 152545 371359
rect 152445 371309 152545 371325
rect 152721 371359 152821 371397
rect 152721 371325 152737 371359
rect 152805 371325 152821 371359
rect 152721 371309 152821 371325
rect 152997 371359 153097 371397
rect 152997 371325 153013 371359
rect 153081 371325 153097 371359
rect 152997 371309 153097 371325
rect 153273 371359 153373 371397
rect 153273 371325 153289 371359
rect 153357 371325 153373 371359
rect 153273 371309 153373 371325
rect 153549 371359 153649 371397
rect 153549 371325 153565 371359
rect 153633 371325 153649 371359
rect 153549 371309 153649 371325
rect 153825 371359 153925 371397
rect 153825 371325 153841 371359
rect 153909 371325 153925 371359
rect 153825 371309 153925 371325
rect 154101 371359 154201 371397
rect 154101 371325 154117 371359
rect 154185 371325 154201 371359
rect 154101 371309 154201 371325
rect 154377 371359 154477 371397
rect 154377 371325 154393 371359
rect 154461 371325 154477 371359
rect 154377 371309 154477 371325
rect 154653 371359 154753 371397
rect 154653 371325 154669 371359
rect 154737 371325 154753 371359
rect 154653 371309 154753 371325
rect 154929 371359 155029 371397
rect 154929 371325 154945 371359
rect 155013 371325 155029 371359
rect 154929 371309 155029 371325
rect 155205 371359 155305 371397
rect 155205 371325 155221 371359
rect 155289 371325 155305 371359
rect 155205 371309 155305 371325
rect 155481 371359 155581 371397
rect 155481 371325 155497 371359
rect 155565 371325 155581 371359
rect 155481 371309 155581 371325
rect 155757 371359 155857 371397
rect 155757 371325 155773 371359
rect 155841 371325 155857 371359
rect 155757 371309 155857 371325
rect 156033 371359 156133 371397
rect 156033 371325 156049 371359
rect 156117 371325 156133 371359
rect 156033 371309 156133 371325
rect 156309 371359 156409 371397
rect 156309 371325 156325 371359
rect 156393 371325 156409 371359
rect 156309 371309 156409 371325
rect 156585 371359 156685 371397
rect 156585 371325 156601 371359
rect 156669 371325 156685 371359
rect 156585 371309 156685 371325
rect 156861 371359 156961 371397
rect 156861 371325 156877 371359
rect 156945 371325 156961 371359
rect 156861 371309 156961 371325
rect 157137 371359 157237 371397
rect 157137 371325 157153 371359
rect 157221 371325 157237 371359
rect 157137 371309 157237 371325
rect 418887 371843 418987 371859
rect 418887 371809 418903 371843
rect 418971 371809 418987 371843
rect 418887 371771 418987 371809
rect 419163 371843 419263 371859
rect 419163 371809 419179 371843
rect 419247 371809 419263 371843
rect 419163 371771 419263 371809
rect 419439 371843 419539 371859
rect 419439 371809 419455 371843
rect 419523 371809 419539 371843
rect 419439 371771 419539 371809
rect 419715 371843 419815 371859
rect 419715 371809 419731 371843
rect 419799 371809 419815 371843
rect 419715 371771 419815 371809
rect 419991 371843 420091 371859
rect 419991 371809 420007 371843
rect 420075 371809 420091 371843
rect 419991 371771 420091 371809
rect 420267 371843 420367 371859
rect 420267 371809 420283 371843
rect 420351 371809 420367 371843
rect 420267 371771 420367 371809
rect 420543 371843 420643 371859
rect 420543 371809 420559 371843
rect 420627 371809 420643 371843
rect 420543 371771 420643 371809
rect 420819 371843 420919 371859
rect 420819 371809 420835 371843
rect 420903 371809 420919 371843
rect 420819 371771 420919 371809
rect 421095 371843 421195 371859
rect 421095 371809 421111 371843
rect 421179 371809 421195 371843
rect 421095 371771 421195 371809
rect 421371 371843 421471 371859
rect 421371 371809 421387 371843
rect 421455 371809 421471 371843
rect 421371 371771 421471 371809
rect 418887 371649 418987 371687
rect 418887 371615 418903 371649
rect 418971 371615 418987 371649
rect 418887 371599 418987 371615
rect 419163 371649 419263 371687
rect 419163 371615 419179 371649
rect 419247 371615 419263 371649
rect 419163 371599 419263 371615
rect 419439 371649 419539 371687
rect 419439 371615 419455 371649
rect 419523 371615 419539 371649
rect 419439 371599 419539 371615
rect 419715 371649 419815 371687
rect 419715 371615 419731 371649
rect 419799 371615 419815 371649
rect 419715 371599 419815 371615
rect 419991 371649 420091 371687
rect 419991 371615 420007 371649
rect 420075 371615 420091 371649
rect 419991 371599 420091 371615
rect 420267 371649 420367 371687
rect 420267 371615 420283 371649
rect 420351 371615 420367 371649
rect 420267 371599 420367 371615
rect 420543 371649 420643 371687
rect 420543 371615 420559 371649
rect 420627 371615 420643 371649
rect 420543 371599 420643 371615
rect 420819 371649 420919 371687
rect 420819 371615 420835 371649
rect 420903 371615 420919 371649
rect 420819 371599 420919 371615
rect 421095 371649 421195 371687
rect 421095 371615 421111 371649
rect 421179 371615 421195 371649
rect 421095 371599 421195 371615
rect 421371 371649 421471 371687
rect 421371 371615 421387 371649
rect 421455 371615 421471 371649
rect 421371 371599 421471 371615
rect 508886 371515 508986 371531
rect 508886 371481 508902 371515
rect 508970 371481 508986 371515
rect 508886 371443 508986 371481
rect 509162 371515 509262 371531
rect 509162 371481 509178 371515
rect 509246 371481 509262 371515
rect 509162 371443 509262 371481
rect 509438 371515 509538 371531
rect 509438 371481 509454 371515
rect 509522 371481 509538 371515
rect 509438 371443 509538 371481
rect 509714 371515 509814 371531
rect 509714 371481 509730 371515
rect 509798 371481 509814 371515
rect 509714 371443 509814 371481
rect 509990 371515 510090 371531
rect 509990 371481 510006 371515
rect 510074 371481 510090 371515
rect 509990 371443 510090 371481
rect 508886 371321 508986 371359
rect 508886 371287 508902 371321
rect 508970 371287 508986 371321
rect 508886 371271 508986 371287
rect 509162 371321 509262 371359
rect 509162 371287 509178 371321
rect 509246 371287 509262 371321
rect 509162 371271 509262 371287
rect 509438 371321 509538 371359
rect 509438 371287 509454 371321
rect 509522 371287 509538 371321
rect 509438 371271 509538 371287
rect 509714 371321 509814 371359
rect 509714 371287 509730 371321
rect 509798 371287 509814 371321
rect 509714 371271 509814 371287
rect 509990 371321 510090 371359
rect 509990 371287 510006 371321
rect 510074 371287 510090 371321
rect 509990 371271 510090 371287
rect 232694 370957 232794 370973
rect 232694 370923 232710 370957
rect 232778 370923 232794 370957
rect 232694 370885 232794 370923
rect 232970 370957 233070 370973
rect 232970 370923 232986 370957
rect 233054 370923 233070 370957
rect 232970 370885 233070 370923
rect 233246 370957 233346 370973
rect 233246 370923 233262 370957
rect 233330 370923 233346 370957
rect 233246 370885 233346 370923
rect 233522 370957 233622 370973
rect 233522 370923 233538 370957
rect 233606 370923 233622 370957
rect 233522 370885 233622 370923
rect 233798 370957 233898 370973
rect 233798 370923 233814 370957
rect 233882 370923 233898 370957
rect 233798 370885 233898 370923
rect 234074 370957 234174 370973
rect 234074 370923 234090 370957
rect 234158 370923 234174 370957
rect 234074 370885 234174 370923
rect 234350 370957 234450 370973
rect 234350 370923 234366 370957
rect 234434 370923 234450 370957
rect 234350 370885 234450 370923
rect 234626 370957 234726 370973
rect 234626 370923 234642 370957
rect 234710 370923 234726 370957
rect 234626 370885 234726 370923
rect 234902 370957 235002 370973
rect 234902 370923 234918 370957
rect 234986 370923 235002 370957
rect 234902 370885 235002 370923
rect 235178 370957 235278 370973
rect 235178 370923 235194 370957
rect 235262 370923 235278 370957
rect 235178 370885 235278 370923
rect 235454 370957 235554 370973
rect 235454 370923 235470 370957
rect 235538 370923 235554 370957
rect 235454 370885 235554 370923
rect 235730 370957 235830 370973
rect 235730 370923 235746 370957
rect 235814 370923 235830 370957
rect 235730 370885 235830 370923
rect 236006 370957 236106 370973
rect 236006 370923 236022 370957
rect 236090 370923 236106 370957
rect 236006 370885 236106 370923
rect 236282 370957 236382 370973
rect 236282 370923 236298 370957
rect 236366 370923 236382 370957
rect 236282 370885 236382 370923
rect 236558 370957 236658 370973
rect 236558 370923 236574 370957
rect 236642 370923 236658 370957
rect 236558 370885 236658 370923
rect 236834 370957 236934 370973
rect 236834 370923 236850 370957
rect 236918 370923 236934 370957
rect 236834 370885 236934 370923
rect 237110 370957 237210 370973
rect 237110 370923 237126 370957
rect 237194 370923 237210 370957
rect 237110 370885 237210 370923
rect 237386 370957 237486 370973
rect 237386 370923 237402 370957
rect 237470 370923 237486 370957
rect 237386 370885 237486 370923
rect 237662 370957 237762 370973
rect 237662 370923 237678 370957
rect 237746 370923 237762 370957
rect 237662 370885 237762 370923
rect 237938 370957 238038 370973
rect 237938 370923 237954 370957
rect 238022 370923 238038 370957
rect 237938 370885 238038 370923
rect 238214 370957 238314 370973
rect 238214 370923 238230 370957
rect 238298 370923 238314 370957
rect 238214 370885 238314 370923
rect 238490 370957 238590 370973
rect 238490 370923 238506 370957
rect 238574 370923 238590 370957
rect 238490 370885 238590 370923
rect 238766 370957 238866 370973
rect 238766 370923 238782 370957
rect 238850 370923 238866 370957
rect 238766 370885 238866 370923
rect 239042 370957 239142 370973
rect 239042 370923 239058 370957
rect 239126 370923 239142 370957
rect 239042 370885 239142 370923
rect 239318 370957 239418 370973
rect 239318 370923 239334 370957
rect 239402 370923 239418 370957
rect 239318 370885 239418 370923
rect 239594 370957 239694 370973
rect 239594 370923 239610 370957
rect 239678 370923 239694 370957
rect 239594 370885 239694 370923
rect 239870 370957 239970 370973
rect 239870 370923 239886 370957
rect 239954 370923 239970 370957
rect 239870 370885 239970 370923
rect 240146 370957 240246 370973
rect 240146 370923 240162 370957
rect 240230 370923 240246 370957
rect 240146 370885 240246 370923
rect 240422 370957 240522 370973
rect 240422 370923 240438 370957
rect 240506 370923 240522 370957
rect 240422 370885 240522 370923
rect 240698 370957 240798 370973
rect 240698 370923 240714 370957
rect 240782 370923 240798 370957
rect 240698 370885 240798 370923
rect 240974 370957 241074 370973
rect 240974 370923 240990 370957
rect 241058 370923 241074 370957
rect 240974 370885 241074 370923
rect 241250 370957 241350 370973
rect 241250 370923 241266 370957
rect 241334 370923 241350 370957
rect 241250 370885 241350 370923
rect 241526 370957 241626 370973
rect 241526 370923 241542 370957
rect 241610 370923 241626 370957
rect 241526 370885 241626 370923
rect 241802 370957 241902 370973
rect 241802 370923 241818 370957
rect 241886 370923 241902 370957
rect 241802 370885 241902 370923
rect 242078 370957 242178 370973
rect 242078 370923 242094 370957
rect 242162 370923 242178 370957
rect 242078 370885 242178 370923
rect 242354 370957 242454 370973
rect 242354 370923 242370 370957
rect 242438 370923 242454 370957
rect 242354 370885 242454 370923
rect 242630 370957 242730 370973
rect 242630 370923 242646 370957
rect 242714 370923 242730 370957
rect 242630 370885 242730 370923
rect 242906 370957 243006 370973
rect 242906 370923 242922 370957
rect 242990 370923 243006 370957
rect 242906 370885 243006 370923
rect 243182 370957 243282 370973
rect 243182 370923 243198 370957
rect 243266 370923 243282 370957
rect 243182 370885 243282 370923
rect 243458 370957 243558 370973
rect 243458 370923 243474 370957
rect 243542 370923 243558 370957
rect 243458 370885 243558 370923
rect 243734 370957 243834 370973
rect 243734 370923 243750 370957
rect 243818 370923 243834 370957
rect 243734 370885 243834 370923
rect 244010 370957 244110 370973
rect 244010 370923 244026 370957
rect 244094 370923 244110 370957
rect 244010 370885 244110 370923
rect 244286 370957 244386 370973
rect 244286 370923 244302 370957
rect 244370 370923 244386 370957
rect 244286 370885 244386 370923
rect 244562 370957 244662 370973
rect 244562 370923 244578 370957
rect 244646 370923 244662 370957
rect 244562 370885 244662 370923
rect 244838 370957 244938 370973
rect 244838 370923 244854 370957
rect 244922 370923 244938 370957
rect 244838 370885 244938 370923
rect 245114 370957 245214 370973
rect 245114 370923 245130 370957
rect 245198 370923 245214 370957
rect 245114 370885 245214 370923
rect 245390 370957 245490 370973
rect 245390 370923 245406 370957
rect 245474 370923 245490 370957
rect 245390 370885 245490 370923
rect 245666 370957 245766 370973
rect 245666 370923 245682 370957
rect 245750 370923 245766 370957
rect 245666 370885 245766 370923
rect 245942 370957 246042 370973
rect 245942 370923 245958 370957
rect 246026 370923 246042 370957
rect 245942 370885 246042 370923
rect 246218 370957 246318 370973
rect 246218 370923 246234 370957
rect 246302 370923 246318 370957
rect 246218 370885 246318 370923
rect 246494 370957 246594 370973
rect 246494 370923 246510 370957
rect 246578 370923 246594 370957
rect 246494 370885 246594 370923
rect 232694 370763 232794 370801
rect 232694 370729 232710 370763
rect 232778 370729 232794 370763
rect 232694 370713 232794 370729
rect 232970 370763 233070 370801
rect 232970 370729 232986 370763
rect 233054 370729 233070 370763
rect 232970 370713 233070 370729
rect 233246 370763 233346 370801
rect 233246 370729 233262 370763
rect 233330 370729 233346 370763
rect 233246 370713 233346 370729
rect 233522 370763 233622 370801
rect 233522 370729 233538 370763
rect 233606 370729 233622 370763
rect 233522 370713 233622 370729
rect 233798 370763 233898 370801
rect 233798 370729 233814 370763
rect 233882 370729 233898 370763
rect 233798 370713 233898 370729
rect 234074 370763 234174 370801
rect 234074 370729 234090 370763
rect 234158 370729 234174 370763
rect 234074 370713 234174 370729
rect 234350 370763 234450 370801
rect 234350 370729 234366 370763
rect 234434 370729 234450 370763
rect 234350 370713 234450 370729
rect 234626 370763 234726 370801
rect 234626 370729 234642 370763
rect 234710 370729 234726 370763
rect 234626 370713 234726 370729
rect 234902 370763 235002 370801
rect 234902 370729 234918 370763
rect 234986 370729 235002 370763
rect 234902 370713 235002 370729
rect 235178 370763 235278 370801
rect 235178 370729 235194 370763
rect 235262 370729 235278 370763
rect 235178 370713 235278 370729
rect 235454 370763 235554 370801
rect 235454 370729 235470 370763
rect 235538 370729 235554 370763
rect 235454 370713 235554 370729
rect 235730 370763 235830 370801
rect 235730 370729 235746 370763
rect 235814 370729 235830 370763
rect 235730 370713 235830 370729
rect 236006 370763 236106 370801
rect 236006 370729 236022 370763
rect 236090 370729 236106 370763
rect 236006 370713 236106 370729
rect 236282 370763 236382 370801
rect 236282 370729 236298 370763
rect 236366 370729 236382 370763
rect 236282 370713 236382 370729
rect 236558 370763 236658 370801
rect 236558 370729 236574 370763
rect 236642 370729 236658 370763
rect 236558 370713 236658 370729
rect 236834 370763 236934 370801
rect 236834 370729 236850 370763
rect 236918 370729 236934 370763
rect 236834 370713 236934 370729
rect 237110 370763 237210 370801
rect 237110 370729 237126 370763
rect 237194 370729 237210 370763
rect 237110 370713 237210 370729
rect 237386 370763 237486 370801
rect 237386 370729 237402 370763
rect 237470 370729 237486 370763
rect 237386 370713 237486 370729
rect 237662 370763 237762 370801
rect 237662 370729 237678 370763
rect 237746 370729 237762 370763
rect 237662 370713 237762 370729
rect 237938 370763 238038 370801
rect 237938 370729 237954 370763
rect 238022 370729 238038 370763
rect 237938 370713 238038 370729
rect 238214 370763 238314 370801
rect 238214 370729 238230 370763
rect 238298 370729 238314 370763
rect 238214 370713 238314 370729
rect 238490 370763 238590 370801
rect 238490 370729 238506 370763
rect 238574 370729 238590 370763
rect 238490 370713 238590 370729
rect 238766 370763 238866 370801
rect 238766 370729 238782 370763
rect 238850 370729 238866 370763
rect 238766 370713 238866 370729
rect 239042 370763 239142 370801
rect 239042 370729 239058 370763
rect 239126 370729 239142 370763
rect 239042 370713 239142 370729
rect 239318 370763 239418 370801
rect 239318 370729 239334 370763
rect 239402 370729 239418 370763
rect 239318 370713 239418 370729
rect 239594 370763 239694 370801
rect 239594 370729 239610 370763
rect 239678 370729 239694 370763
rect 239594 370713 239694 370729
rect 239870 370763 239970 370801
rect 239870 370729 239886 370763
rect 239954 370729 239970 370763
rect 239870 370713 239970 370729
rect 240146 370763 240246 370801
rect 240146 370729 240162 370763
rect 240230 370729 240246 370763
rect 240146 370713 240246 370729
rect 240422 370763 240522 370801
rect 240422 370729 240438 370763
rect 240506 370729 240522 370763
rect 240422 370713 240522 370729
rect 240698 370763 240798 370801
rect 240698 370729 240714 370763
rect 240782 370729 240798 370763
rect 240698 370713 240798 370729
rect 240974 370763 241074 370801
rect 240974 370729 240990 370763
rect 241058 370729 241074 370763
rect 240974 370713 241074 370729
rect 241250 370763 241350 370801
rect 241250 370729 241266 370763
rect 241334 370729 241350 370763
rect 241250 370713 241350 370729
rect 241526 370763 241626 370801
rect 241526 370729 241542 370763
rect 241610 370729 241626 370763
rect 241526 370713 241626 370729
rect 241802 370763 241902 370801
rect 241802 370729 241818 370763
rect 241886 370729 241902 370763
rect 241802 370713 241902 370729
rect 242078 370763 242178 370801
rect 242078 370729 242094 370763
rect 242162 370729 242178 370763
rect 242078 370713 242178 370729
rect 242354 370763 242454 370801
rect 242354 370729 242370 370763
rect 242438 370729 242454 370763
rect 242354 370713 242454 370729
rect 242630 370763 242730 370801
rect 242630 370729 242646 370763
rect 242714 370729 242730 370763
rect 242630 370713 242730 370729
rect 242906 370763 243006 370801
rect 242906 370729 242922 370763
rect 242990 370729 243006 370763
rect 242906 370713 243006 370729
rect 243182 370763 243282 370801
rect 243182 370729 243198 370763
rect 243266 370729 243282 370763
rect 243182 370713 243282 370729
rect 243458 370763 243558 370801
rect 243458 370729 243474 370763
rect 243542 370729 243558 370763
rect 243458 370713 243558 370729
rect 243734 370763 243834 370801
rect 243734 370729 243750 370763
rect 243818 370729 243834 370763
rect 243734 370713 243834 370729
rect 244010 370763 244110 370801
rect 244010 370729 244026 370763
rect 244094 370729 244110 370763
rect 244010 370713 244110 370729
rect 244286 370763 244386 370801
rect 244286 370729 244302 370763
rect 244370 370729 244386 370763
rect 244286 370713 244386 370729
rect 244562 370763 244662 370801
rect 244562 370729 244578 370763
rect 244646 370729 244662 370763
rect 244562 370713 244662 370729
rect 244838 370763 244938 370801
rect 244838 370729 244854 370763
rect 244922 370729 244938 370763
rect 244838 370713 244938 370729
rect 245114 370763 245214 370801
rect 245114 370729 245130 370763
rect 245198 370729 245214 370763
rect 245114 370713 245214 370729
rect 245390 370763 245490 370801
rect 245390 370729 245406 370763
rect 245474 370729 245490 370763
rect 245390 370713 245490 370729
rect 245666 370763 245766 370801
rect 245666 370729 245682 370763
rect 245750 370729 245766 370763
rect 245666 370713 245766 370729
rect 245942 370763 246042 370801
rect 245942 370729 245958 370763
rect 246026 370729 246042 370763
rect 245942 370713 246042 370729
rect 246218 370763 246318 370801
rect 246218 370729 246234 370763
rect 246302 370729 246318 370763
rect 246218 370713 246318 370729
rect 246494 370763 246594 370801
rect 246494 370729 246510 370763
rect 246578 370729 246594 370763
rect 246494 370713 246594 370729
rect 58886 251515 58986 251531
rect 58886 251481 58902 251515
rect 58970 251481 58986 251515
rect 58886 251443 58986 251481
rect 59162 251515 59262 251531
rect 59162 251481 59178 251515
rect 59246 251481 59262 251515
rect 59162 251443 59262 251481
rect 59438 251515 59538 251531
rect 59438 251481 59454 251515
rect 59522 251481 59538 251515
rect 59438 251443 59538 251481
rect 59714 251515 59814 251531
rect 59714 251481 59730 251515
rect 59798 251481 59814 251515
rect 59714 251443 59814 251481
rect 59990 251515 60090 251531
rect 59990 251481 60006 251515
rect 60074 251481 60090 251515
rect 59990 251443 60090 251481
rect 58886 251321 58986 251359
rect 58886 251287 58902 251321
rect 58970 251287 58986 251321
rect 58886 251271 58986 251287
rect 59162 251321 59262 251359
rect 59162 251287 59178 251321
rect 59246 251287 59262 251321
rect 59162 251271 59262 251287
rect 59438 251321 59538 251359
rect 59438 251287 59454 251321
rect 59522 251287 59538 251321
rect 59438 251271 59538 251287
rect 59714 251321 59814 251359
rect 59714 251287 59730 251321
rect 59798 251287 59814 251321
rect 59714 251271 59814 251287
rect 59990 251321 60090 251359
rect 59990 251287 60006 251321
rect 60074 251287 60090 251321
rect 59990 251271 60090 251287
rect 148011 251639 148111 251655
rect 148011 251605 148027 251639
rect 148095 251605 148111 251639
rect 148011 251567 148111 251605
rect 148287 251639 148387 251655
rect 148287 251605 148303 251639
rect 148371 251605 148387 251639
rect 148287 251567 148387 251605
rect 148563 251639 148663 251655
rect 148563 251605 148579 251639
rect 148647 251605 148663 251639
rect 148563 251567 148663 251605
rect 148839 251639 148939 251655
rect 148839 251605 148855 251639
rect 148923 251605 148939 251639
rect 148839 251567 148939 251605
rect 149115 251639 149215 251655
rect 149115 251605 149131 251639
rect 149199 251605 149215 251639
rect 149115 251567 149215 251605
rect 149391 251639 149491 251655
rect 149391 251605 149407 251639
rect 149475 251605 149491 251639
rect 149391 251567 149491 251605
rect 149667 251639 149767 251655
rect 149667 251605 149683 251639
rect 149751 251605 149767 251639
rect 149667 251567 149767 251605
rect 149943 251639 150043 251655
rect 149943 251605 149959 251639
rect 150027 251605 150043 251639
rect 149943 251567 150043 251605
rect 150219 251639 150319 251655
rect 150219 251605 150235 251639
rect 150303 251605 150319 251639
rect 150219 251567 150319 251605
rect 150495 251639 150595 251655
rect 150495 251605 150511 251639
rect 150579 251605 150595 251639
rect 150495 251567 150595 251605
rect 148011 251445 148111 251483
rect 148011 251411 148027 251445
rect 148095 251411 148111 251445
rect 148011 251395 148111 251411
rect 148287 251445 148387 251483
rect 148287 251411 148303 251445
rect 148371 251411 148387 251445
rect 148287 251395 148387 251411
rect 148563 251445 148663 251483
rect 148563 251411 148579 251445
rect 148647 251411 148663 251445
rect 148563 251395 148663 251411
rect 148839 251445 148939 251483
rect 148839 251411 148855 251445
rect 148923 251411 148939 251445
rect 148839 251395 148939 251411
rect 149115 251445 149215 251483
rect 149115 251411 149131 251445
rect 149199 251411 149215 251445
rect 149115 251395 149215 251411
rect 149391 251445 149491 251483
rect 149391 251411 149407 251445
rect 149475 251411 149491 251445
rect 149391 251395 149491 251411
rect 149667 251445 149767 251483
rect 149667 251411 149683 251445
rect 149751 251411 149767 251445
rect 149667 251395 149767 251411
rect 149943 251445 150043 251483
rect 149943 251411 149959 251445
rect 150027 251411 150043 251445
rect 149943 251395 150043 251411
rect 150219 251445 150319 251483
rect 150219 251411 150235 251445
rect 150303 251411 150319 251445
rect 150219 251395 150319 251411
rect 150495 251445 150595 251483
rect 150495 251411 150511 251445
rect 150579 251411 150595 251445
rect 150495 251395 150595 251411
rect 234255 251839 234355 251855
rect 234255 251805 234271 251839
rect 234339 251805 234355 251839
rect 234255 251767 234355 251805
rect 234531 251839 234631 251855
rect 234531 251805 234547 251839
rect 234615 251805 234631 251839
rect 234531 251767 234631 251805
rect 234807 251839 234907 251855
rect 234807 251805 234823 251839
rect 234891 251805 234907 251839
rect 234807 251767 234907 251805
rect 235083 251839 235183 251855
rect 235083 251805 235099 251839
rect 235167 251805 235183 251839
rect 235083 251767 235183 251805
rect 235359 251839 235459 251855
rect 235359 251805 235375 251839
rect 235443 251805 235459 251839
rect 235359 251767 235459 251805
rect 235635 251839 235735 251855
rect 235635 251805 235651 251839
rect 235719 251805 235735 251839
rect 235635 251767 235735 251805
rect 235911 251839 236011 251855
rect 235911 251805 235927 251839
rect 235995 251805 236011 251839
rect 235911 251767 236011 251805
rect 236187 251839 236287 251855
rect 236187 251805 236203 251839
rect 236271 251805 236287 251839
rect 236187 251767 236287 251805
rect 236463 251839 236563 251855
rect 236463 251805 236479 251839
rect 236547 251805 236563 251839
rect 236463 251767 236563 251805
rect 236739 251839 236839 251855
rect 236739 251805 236755 251839
rect 236823 251805 236839 251839
rect 236739 251767 236839 251805
rect 237015 251839 237115 251855
rect 237015 251805 237031 251839
rect 237099 251805 237115 251839
rect 237015 251767 237115 251805
rect 237291 251839 237391 251855
rect 237291 251805 237307 251839
rect 237375 251805 237391 251839
rect 237291 251767 237391 251805
rect 237567 251839 237667 251855
rect 237567 251805 237583 251839
rect 237651 251805 237667 251839
rect 237567 251767 237667 251805
rect 237843 251839 237943 251855
rect 237843 251805 237859 251839
rect 237927 251805 237943 251839
rect 237843 251767 237943 251805
rect 238119 251839 238219 251855
rect 238119 251805 238135 251839
rect 238203 251805 238219 251839
rect 238119 251767 238219 251805
rect 238395 251839 238495 251855
rect 238395 251805 238411 251839
rect 238479 251805 238495 251839
rect 238395 251767 238495 251805
rect 238671 251839 238771 251855
rect 238671 251805 238687 251839
rect 238755 251805 238771 251839
rect 238671 251767 238771 251805
rect 238947 251839 239047 251855
rect 238947 251805 238963 251839
rect 239031 251805 239047 251839
rect 238947 251767 239047 251805
rect 239223 251839 239323 251855
rect 239223 251805 239239 251839
rect 239307 251805 239323 251839
rect 239223 251767 239323 251805
rect 239499 251839 239599 251855
rect 239499 251805 239515 251839
rect 239583 251805 239599 251839
rect 239499 251767 239599 251805
rect 239775 251839 239875 251855
rect 239775 251805 239791 251839
rect 239859 251805 239875 251839
rect 239775 251767 239875 251805
rect 240051 251839 240151 251855
rect 240051 251805 240067 251839
rect 240135 251805 240151 251839
rect 240051 251767 240151 251805
rect 240327 251839 240427 251855
rect 240327 251805 240343 251839
rect 240411 251805 240427 251839
rect 240327 251767 240427 251805
rect 240603 251839 240703 251855
rect 240603 251805 240619 251839
rect 240687 251805 240703 251839
rect 240603 251767 240703 251805
rect 240879 251839 240979 251855
rect 240879 251805 240895 251839
rect 240963 251805 240979 251839
rect 240879 251767 240979 251805
rect 241155 251839 241255 251855
rect 241155 251805 241171 251839
rect 241239 251805 241255 251839
rect 241155 251767 241255 251805
rect 241431 251839 241531 251855
rect 241431 251805 241447 251839
rect 241515 251805 241531 251839
rect 241431 251767 241531 251805
rect 241707 251839 241807 251855
rect 241707 251805 241723 251839
rect 241791 251805 241807 251839
rect 241707 251767 241807 251805
rect 241983 251839 242083 251855
rect 241983 251805 241999 251839
rect 242067 251805 242083 251839
rect 241983 251767 242083 251805
rect 242259 251839 242359 251855
rect 242259 251805 242275 251839
rect 242343 251805 242359 251839
rect 242259 251767 242359 251805
rect 242535 251839 242635 251855
rect 242535 251805 242551 251839
rect 242619 251805 242635 251839
rect 242535 251767 242635 251805
rect 242811 251839 242911 251855
rect 242811 251805 242827 251839
rect 242895 251805 242911 251839
rect 242811 251767 242911 251805
rect 243087 251839 243187 251855
rect 243087 251805 243103 251839
rect 243171 251805 243187 251839
rect 243087 251767 243187 251805
rect 243363 251839 243463 251855
rect 243363 251805 243379 251839
rect 243447 251805 243463 251839
rect 243363 251767 243463 251805
rect 243639 251839 243739 251855
rect 243639 251805 243655 251839
rect 243723 251805 243739 251839
rect 243639 251767 243739 251805
rect 243915 251839 244015 251855
rect 243915 251805 243931 251839
rect 243999 251805 244015 251839
rect 243915 251767 244015 251805
rect 244191 251839 244291 251855
rect 244191 251805 244207 251839
rect 244275 251805 244291 251839
rect 244191 251767 244291 251805
rect 244467 251839 244567 251855
rect 244467 251805 244483 251839
rect 244551 251805 244567 251839
rect 244467 251767 244567 251805
rect 244743 251839 244843 251855
rect 244743 251805 244759 251839
rect 244827 251805 244843 251839
rect 244743 251767 244843 251805
rect 245019 251839 245119 251855
rect 245019 251805 245035 251839
rect 245103 251805 245119 251839
rect 245019 251767 245119 251805
rect 245295 251839 245395 251855
rect 245295 251805 245311 251839
rect 245379 251805 245395 251839
rect 245295 251767 245395 251805
rect 245571 251839 245671 251855
rect 245571 251805 245587 251839
rect 245655 251805 245671 251839
rect 245571 251767 245671 251805
rect 245847 251839 245947 251855
rect 245847 251805 245863 251839
rect 245931 251805 245947 251839
rect 245847 251767 245947 251805
rect 246123 251839 246223 251855
rect 246123 251805 246139 251839
rect 246207 251805 246223 251839
rect 246123 251767 246223 251805
rect 246399 251839 246499 251855
rect 246399 251805 246415 251839
rect 246483 251805 246499 251839
rect 246399 251767 246499 251805
rect 246675 251839 246775 251855
rect 246675 251805 246691 251839
rect 246759 251805 246775 251839
rect 246675 251767 246775 251805
rect 246951 251839 247051 251855
rect 246951 251805 246967 251839
rect 247035 251805 247051 251839
rect 246951 251767 247051 251805
rect 247227 251839 247327 251855
rect 247227 251805 247243 251839
rect 247311 251805 247327 251839
rect 247227 251767 247327 251805
rect 247503 251839 247603 251855
rect 247503 251805 247519 251839
rect 247587 251805 247603 251839
rect 247503 251767 247603 251805
rect 247779 251839 247879 251855
rect 247779 251805 247795 251839
rect 247863 251805 247879 251839
rect 247779 251767 247879 251805
rect 248055 251839 248155 251855
rect 248055 251805 248071 251839
rect 248139 251805 248155 251839
rect 248055 251767 248155 251805
rect 234255 251645 234355 251683
rect 234255 251611 234271 251645
rect 234339 251611 234355 251645
rect 234255 251595 234355 251611
rect 234531 251645 234631 251683
rect 234531 251611 234547 251645
rect 234615 251611 234631 251645
rect 234531 251595 234631 251611
rect 234807 251645 234907 251683
rect 234807 251611 234823 251645
rect 234891 251611 234907 251645
rect 234807 251595 234907 251611
rect 235083 251645 235183 251683
rect 235083 251611 235099 251645
rect 235167 251611 235183 251645
rect 235083 251595 235183 251611
rect 235359 251645 235459 251683
rect 235359 251611 235375 251645
rect 235443 251611 235459 251645
rect 235359 251595 235459 251611
rect 235635 251645 235735 251683
rect 235635 251611 235651 251645
rect 235719 251611 235735 251645
rect 235635 251595 235735 251611
rect 235911 251645 236011 251683
rect 235911 251611 235927 251645
rect 235995 251611 236011 251645
rect 235911 251595 236011 251611
rect 236187 251645 236287 251683
rect 236187 251611 236203 251645
rect 236271 251611 236287 251645
rect 236187 251595 236287 251611
rect 236463 251645 236563 251683
rect 236463 251611 236479 251645
rect 236547 251611 236563 251645
rect 236463 251595 236563 251611
rect 236739 251645 236839 251683
rect 236739 251611 236755 251645
rect 236823 251611 236839 251645
rect 236739 251595 236839 251611
rect 237015 251645 237115 251683
rect 237015 251611 237031 251645
rect 237099 251611 237115 251645
rect 237015 251595 237115 251611
rect 237291 251645 237391 251683
rect 237291 251611 237307 251645
rect 237375 251611 237391 251645
rect 237291 251595 237391 251611
rect 237567 251645 237667 251683
rect 237567 251611 237583 251645
rect 237651 251611 237667 251645
rect 237567 251595 237667 251611
rect 237843 251645 237943 251683
rect 237843 251611 237859 251645
rect 237927 251611 237943 251645
rect 237843 251595 237943 251611
rect 238119 251645 238219 251683
rect 238119 251611 238135 251645
rect 238203 251611 238219 251645
rect 238119 251595 238219 251611
rect 238395 251645 238495 251683
rect 238395 251611 238411 251645
rect 238479 251611 238495 251645
rect 238395 251595 238495 251611
rect 238671 251645 238771 251683
rect 238671 251611 238687 251645
rect 238755 251611 238771 251645
rect 238671 251595 238771 251611
rect 238947 251645 239047 251683
rect 238947 251611 238963 251645
rect 239031 251611 239047 251645
rect 238947 251595 239047 251611
rect 239223 251645 239323 251683
rect 239223 251611 239239 251645
rect 239307 251611 239323 251645
rect 239223 251595 239323 251611
rect 239499 251645 239599 251683
rect 239499 251611 239515 251645
rect 239583 251611 239599 251645
rect 239499 251595 239599 251611
rect 239775 251645 239875 251683
rect 239775 251611 239791 251645
rect 239859 251611 239875 251645
rect 239775 251595 239875 251611
rect 240051 251645 240151 251683
rect 240051 251611 240067 251645
rect 240135 251611 240151 251645
rect 240051 251595 240151 251611
rect 240327 251645 240427 251683
rect 240327 251611 240343 251645
rect 240411 251611 240427 251645
rect 240327 251595 240427 251611
rect 240603 251645 240703 251683
rect 240603 251611 240619 251645
rect 240687 251611 240703 251645
rect 240603 251595 240703 251611
rect 240879 251645 240979 251683
rect 240879 251611 240895 251645
rect 240963 251611 240979 251645
rect 240879 251595 240979 251611
rect 241155 251645 241255 251683
rect 241155 251611 241171 251645
rect 241239 251611 241255 251645
rect 241155 251595 241255 251611
rect 241431 251645 241531 251683
rect 241431 251611 241447 251645
rect 241515 251611 241531 251645
rect 241431 251595 241531 251611
rect 241707 251645 241807 251683
rect 241707 251611 241723 251645
rect 241791 251611 241807 251645
rect 241707 251595 241807 251611
rect 241983 251645 242083 251683
rect 241983 251611 241999 251645
rect 242067 251611 242083 251645
rect 241983 251595 242083 251611
rect 242259 251645 242359 251683
rect 242259 251611 242275 251645
rect 242343 251611 242359 251645
rect 242259 251595 242359 251611
rect 242535 251645 242635 251683
rect 242535 251611 242551 251645
rect 242619 251611 242635 251645
rect 242535 251595 242635 251611
rect 242811 251645 242911 251683
rect 242811 251611 242827 251645
rect 242895 251611 242911 251645
rect 242811 251595 242911 251611
rect 243087 251645 243187 251683
rect 243087 251611 243103 251645
rect 243171 251611 243187 251645
rect 243087 251595 243187 251611
rect 243363 251645 243463 251683
rect 243363 251611 243379 251645
rect 243447 251611 243463 251645
rect 243363 251595 243463 251611
rect 243639 251645 243739 251683
rect 243639 251611 243655 251645
rect 243723 251611 243739 251645
rect 243639 251595 243739 251611
rect 243915 251645 244015 251683
rect 243915 251611 243931 251645
rect 243999 251611 244015 251645
rect 243915 251595 244015 251611
rect 244191 251645 244291 251683
rect 244191 251611 244207 251645
rect 244275 251611 244291 251645
rect 244191 251595 244291 251611
rect 244467 251645 244567 251683
rect 244467 251611 244483 251645
rect 244551 251611 244567 251645
rect 244467 251595 244567 251611
rect 244743 251645 244843 251683
rect 244743 251611 244759 251645
rect 244827 251611 244843 251645
rect 244743 251595 244843 251611
rect 245019 251645 245119 251683
rect 245019 251611 245035 251645
rect 245103 251611 245119 251645
rect 245019 251595 245119 251611
rect 245295 251645 245395 251683
rect 245295 251611 245311 251645
rect 245379 251611 245395 251645
rect 245295 251595 245395 251611
rect 245571 251645 245671 251683
rect 245571 251611 245587 251645
rect 245655 251611 245671 251645
rect 245571 251595 245671 251611
rect 245847 251645 245947 251683
rect 245847 251611 245863 251645
rect 245931 251611 245947 251645
rect 245847 251595 245947 251611
rect 246123 251645 246223 251683
rect 246123 251611 246139 251645
rect 246207 251611 246223 251645
rect 246123 251595 246223 251611
rect 246399 251645 246499 251683
rect 246399 251611 246415 251645
rect 246483 251611 246499 251645
rect 246399 251595 246499 251611
rect 246675 251645 246775 251683
rect 246675 251611 246691 251645
rect 246759 251611 246775 251645
rect 246675 251595 246775 251611
rect 246951 251645 247051 251683
rect 246951 251611 246967 251645
rect 247035 251611 247051 251645
rect 246951 251595 247051 251611
rect 247227 251645 247327 251683
rect 247227 251611 247243 251645
rect 247311 251611 247327 251645
rect 247227 251595 247327 251611
rect 247503 251645 247603 251683
rect 247503 251611 247519 251645
rect 247587 251611 247603 251645
rect 247503 251595 247603 251611
rect 247779 251645 247879 251683
rect 247779 251611 247795 251645
rect 247863 251611 247879 251645
rect 247779 251595 247879 251611
rect 248055 251645 248155 251683
rect 248055 251611 248071 251645
rect 248139 251611 248155 251645
rect 248055 251595 248155 251611
rect 413337 251553 413437 251569
rect 413337 251519 413353 251553
rect 413421 251519 413437 251553
rect 413337 251481 413437 251519
rect 413613 251553 413713 251569
rect 413613 251519 413629 251553
rect 413697 251519 413713 251553
rect 413613 251481 413713 251519
rect 413889 251553 413989 251569
rect 413889 251519 413905 251553
rect 413973 251519 413989 251553
rect 413889 251481 413989 251519
rect 414165 251553 414265 251569
rect 414165 251519 414181 251553
rect 414249 251519 414265 251553
rect 414165 251481 414265 251519
rect 414441 251553 414541 251569
rect 414441 251519 414457 251553
rect 414525 251519 414541 251553
rect 414441 251481 414541 251519
rect 414717 251553 414817 251569
rect 414717 251519 414733 251553
rect 414801 251519 414817 251553
rect 414717 251481 414817 251519
rect 414993 251553 415093 251569
rect 414993 251519 415009 251553
rect 415077 251519 415093 251553
rect 414993 251481 415093 251519
rect 415269 251553 415369 251569
rect 415269 251519 415285 251553
rect 415353 251519 415369 251553
rect 415269 251481 415369 251519
rect 415545 251553 415645 251569
rect 415545 251519 415561 251553
rect 415629 251519 415645 251553
rect 415545 251481 415645 251519
rect 415821 251553 415921 251569
rect 415821 251519 415837 251553
rect 415905 251519 415921 251553
rect 415821 251481 415921 251519
rect 416097 251553 416197 251569
rect 416097 251519 416113 251553
rect 416181 251519 416197 251553
rect 416097 251481 416197 251519
rect 416373 251553 416473 251569
rect 416373 251519 416389 251553
rect 416457 251519 416473 251553
rect 416373 251481 416473 251519
rect 416649 251553 416749 251569
rect 416649 251519 416665 251553
rect 416733 251519 416749 251553
rect 416649 251481 416749 251519
rect 416925 251553 417025 251569
rect 416925 251519 416941 251553
rect 417009 251519 417025 251553
rect 416925 251481 417025 251519
rect 417201 251553 417301 251569
rect 417201 251519 417217 251553
rect 417285 251519 417301 251553
rect 417201 251481 417301 251519
rect 417477 251553 417577 251569
rect 417477 251519 417493 251553
rect 417561 251519 417577 251553
rect 417477 251481 417577 251519
rect 417753 251553 417853 251569
rect 417753 251519 417769 251553
rect 417837 251519 417853 251553
rect 417753 251481 417853 251519
rect 418029 251553 418129 251569
rect 418029 251519 418045 251553
rect 418113 251519 418129 251553
rect 418029 251481 418129 251519
rect 418305 251553 418405 251569
rect 418305 251519 418321 251553
rect 418389 251519 418405 251553
rect 418305 251481 418405 251519
rect 418581 251553 418681 251569
rect 418581 251519 418597 251553
rect 418665 251519 418681 251553
rect 418581 251481 418681 251519
rect 418857 251553 418957 251569
rect 418857 251519 418873 251553
rect 418941 251519 418957 251553
rect 418857 251481 418957 251519
rect 419133 251553 419233 251569
rect 419133 251519 419149 251553
rect 419217 251519 419233 251553
rect 419133 251481 419233 251519
rect 419409 251553 419509 251569
rect 419409 251519 419425 251553
rect 419493 251519 419509 251553
rect 419409 251481 419509 251519
rect 419685 251553 419785 251569
rect 419685 251519 419701 251553
rect 419769 251519 419785 251553
rect 419685 251481 419785 251519
rect 419961 251553 420061 251569
rect 419961 251519 419977 251553
rect 420045 251519 420061 251553
rect 419961 251481 420061 251519
rect 420237 251553 420337 251569
rect 420237 251519 420253 251553
rect 420321 251519 420337 251553
rect 420237 251481 420337 251519
rect 420513 251553 420613 251569
rect 420513 251519 420529 251553
rect 420597 251519 420613 251553
rect 420513 251481 420613 251519
rect 420789 251553 420889 251569
rect 420789 251519 420805 251553
rect 420873 251519 420889 251553
rect 420789 251481 420889 251519
rect 421065 251553 421165 251569
rect 421065 251519 421081 251553
rect 421149 251519 421165 251553
rect 421065 251481 421165 251519
rect 421341 251553 421441 251569
rect 421341 251519 421357 251553
rect 421425 251519 421441 251553
rect 421341 251481 421441 251519
rect 421617 251553 421717 251569
rect 421617 251519 421633 251553
rect 421701 251519 421717 251553
rect 421617 251481 421717 251519
rect 421893 251553 421993 251569
rect 421893 251519 421909 251553
rect 421977 251519 421993 251553
rect 421893 251481 421993 251519
rect 422169 251553 422269 251569
rect 422169 251519 422185 251553
rect 422253 251519 422269 251553
rect 422169 251481 422269 251519
rect 422445 251553 422545 251569
rect 422445 251519 422461 251553
rect 422529 251519 422545 251553
rect 422445 251481 422545 251519
rect 422721 251553 422821 251569
rect 422721 251519 422737 251553
rect 422805 251519 422821 251553
rect 422721 251481 422821 251519
rect 422997 251553 423097 251569
rect 422997 251519 423013 251553
rect 423081 251519 423097 251553
rect 422997 251481 423097 251519
rect 423273 251553 423373 251569
rect 423273 251519 423289 251553
rect 423357 251519 423373 251553
rect 423273 251481 423373 251519
rect 423549 251553 423649 251569
rect 423549 251519 423565 251553
rect 423633 251519 423649 251553
rect 423549 251481 423649 251519
rect 423825 251553 423925 251569
rect 423825 251519 423841 251553
rect 423909 251519 423925 251553
rect 423825 251481 423925 251519
rect 424101 251553 424201 251569
rect 424101 251519 424117 251553
rect 424185 251519 424201 251553
rect 424101 251481 424201 251519
rect 424377 251553 424477 251569
rect 424377 251519 424393 251553
rect 424461 251519 424477 251553
rect 424377 251481 424477 251519
rect 424653 251553 424753 251569
rect 424653 251519 424669 251553
rect 424737 251519 424753 251553
rect 424653 251481 424753 251519
rect 424929 251553 425029 251569
rect 424929 251519 424945 251553
rect 425013 251519 425029 251553
rect 424929 251481 425029 251519
rect 425205 251553 425305 251569
rect 425205 251519 425221 251553
rect 425289 251519 425305 251553
rect 425205 251481 425305 251519
rect 425481 251553 425581 251569
rect 425481 251519 425497 251553
rect 425565 251519 425581 251553
rect 425481 251481 425581 251519
rect 425757 251553 425857 251569
rect 425757 251519 425773 251553
rect 425841 251519 425857 251553
rect 425757 251481 425857 251519
rect 426033 251553 426133 251569
rect 426033 251519 426049 251553
rect 426117 251519 426133 251553
rect 426033 251481 426133 251519
rect 426309 251553 426409 251569
rect 426309 251519 426325 251553
rect 426393 251519 426409 251553
rect 426309 251481 426409 251519
rect 426585 251553 426685 251569
rect 426585 251519 426601 251553
rect 426669 251519 426685 251553
rect 426585 251481 426685 251519
rect 426861 251553 426961 251569
rect 426861 251519 426877 251553
rect 426945 251519 426961 251553
rect 426861 251481 426961 251519
rect 427137 251553 427237 251569
rect 427137 251519 427153 251553
rect 427221 251519 427237 251553
rect 427137 251481 427237 251519
rect 413337 251359 413437 251397
rect 413337 251325 413353 251359
rect 413421 251325 413437 251359
rect 413337 251309 413437 251325
rect 413613 251359 413713 251397
rect 413613 251325 413629 251359
rect 413697 251325 413713 251359
rect 413613 251309 413713 251325
rect 413889 251359 413989 251397
rect 413889 251325 413905 251359
rect 413973 251325 413989 251359
rect 413889 251309 413989 251325
rect 414165 251359 414265 251397
rect 414165 251325 414181 251359
rect 414249 251325 414265 251359
rect 414165 251309 414265 251325
rect 414441 251359 414541 251397
rect 414441 251325 414457 251359
rect 414525 251325 414541 251359
rect 414441 251309 414541 251325
rect 414717 251359 414817 251397
rect 414717 251325 414733 251359
rect 414801 251325 414817 251359
rect 414717 251309 414817 251325
rect 414993 251359 415093 251397
rect 414993 251325 415009 251359
rect 415077 251325 415093 251359
rect 414993 251309 415093 251325
rect 415269 251359 415369 251397
rect 415269 251325 415285 251359
rect 415353 251325 415369 251359
rect 415269 251309 415369 251325
rect 415545 251359 415645 251397
rect 415545 251325 415561 251359
rect 415629 251325 415645 251359
rect 415545 251309 415645 251325
rect 415821 251359 415921 251397
rect 415821 251325 415837 251359
rect 415905 251325 415921 251359
rect 415821 251309 415921 251325
rect 416097 251359 416197 251397
rect 416097 251325 416113 251359
rect 416181 251325 416197 251359
rect 416097 251309 416197 251325
rect 416373 251359 416473 251397
rect 416373 251325 416389 251359
rect 416457 251325 416473 251359
rect 416373 251309 416473 251325
rect 416649 251359 416749 251397
rect 416649 251325 416665 251359
rect 416733 251325 416749 251359
rect 416649 251309 416749 251325
rect 416925 251359 417025 251397
rect 416925 251325 416941 251359
rect 417009 251325 417025 251359
rect 416925 251309 417025 251325
rect 417201 251359 417301 251397
rect 417201 251325 417217 251359
rect 417285 251325 417301 251359
rect 417201 251309 417301 251325
rect 417477 251359 417577 251397
rect 417477 251325 417493 251359
rect 417561 251325 417577 251359
rect 417477 251309 417577 251325
rect 417753 251359 417853 251397
rect 417753 251325 417769 251359
rect 417837 251325 417853 251359
rect 417753 251309 417853 251325
rect 418029 251359 418129 251397
rect 418029 251325 418045 251359
rect 418113 251325 418129 251359
rect 418029 251309 418129 251325
rect 418305 251359 418405 251397
rect 418305 251325 418321 251359
rect 418389 251325 418405 251359
rect 418305 251309 418405 251325
rect 418581 251359 418681 251397
rect 418581 251325 418597 251359
rect 418665 251325 418681 251359
rect 418581 251309 418681 251325
rect 418857 251359 418957 251397
rect 418857 251325 418873 251359
rect 418941 251325 418957 251359
rect 418857 251309 418957 251325
rect 419133 251359 419233 251397
rect 419133 251325 419149 251359
rect 419217 251325 419233 251359
rect 419133 251309 419233 251325
rect 419409 251359 419509 251397
rect 419409 251325 419425 251359
rect 419493 251325 419509 251359
rect 419409 251309 419509 251325
rect 419685 251359 419785 251397
rect 419685 251325 419701 251359
rect 419769 251325 419785 251359
rect 419685 251309 419785 251325
rect 419961 251359 420061 251397
rect 419961 251325 419977 251359
rect 420045 251325 420061 251359
rect 419961 251309 420061 251325
rect 420237 251359 420337 251397
rect 420237 251325 420253 251359
rect 420321 251325 420337 251359
rect 420237 251309 420337 251325
rect 420513 251359 420613 251397
rect 420513 251325 420529 251359
rect 420597 251325 420613 251359
rect 420513 251309 420613 251325
rect 420789 251359 420889 251397
rect 420789 251325 420805 251359
rect 420873 251325 420889 251359
rect 420789 251309 420889 251325
rect 421065 251359 421165 251397
rect 421065 251325 421081 251359
rect 421149 251325 421165 251359
rect 421065 251309 421165 251325
rect 421341 251359 421441 251397
rect 421341 251325 421357 251359
rect 421425 251325 421441 251359
rect 421341 251309 421441 251325
rect 421617 251359 421717 251397
rect 421617 251325 421633 251359
rect 421701 251325 421717 251359
rect 421617 251309 421717 251325
rect 421893 251359 421993 251397
rect 421893 251325 421909 251359
rect 421977 251325 421993 251359
rect 421893 251309 421993 251325
rect 422169 251359 422269 251397
rect 422169 251325 422185 251359
rect 422253 251325 422269 251359
rect 422169 251309 422269 251325
rect 422445 251359 422545 251397
rect 422445 251325 422461 251359
rect 422529 251325 422545 251359
rect 422445 251309 422545 251325
rect 422721 251359 422821 251397
rect 422721 251325 422737 251359
rect 422805 251325 422821 251359
rect 422721 251309 422821 251325
rect 422997 251359 423097 251397
rect 422997 251325 423013 251359
rect 423081 251325 423097 251359
rect 422997 251309 423097 251325
rect 423273 251359 423373 251397
rect 423273 251325 423289 251359
rect 423357 251325 423373 251359
rect 423273 251309 423373 251325
rect 423549 251359 423649 251397
rect 423549 251325 423565 251359
rect 423633 251325 423649 251359
rect 423549 251309 423649 251325
rect 423825 251359 423925 251397
rect 423825 251325 423841 251359
rect 423909 251325 423925 251359
rect 423825 251309 423925 251325
rect 424101 251359 424201 251397
rect 424101 251325 424117 251359
rect 424185 251325 424201 251359
rect 424101 251309 424201 251325
rect 424377 251359 424477 251397
rect 424377 251325 424393 251359
rect 424461 251325 424477 251359
rect 424377 251309 424477 251325
rect 424653 251359 424753 251397
rect 424653 251325 424669 251359
rect 424737 251325 424753 251359
rect 424653 251309 424753 251325
rect 424929 251359 425029 251397
rect 424929 251325 424945 251359
rect 425013 251325 425029 251359
rect 424929 251309 425029 251325
rect 425205 251359 425305 251397
rect 425205 251325 425221 251359
rect 425289 251325 425305 251359
rect 425205 251309 425305 251325
rect 425481 251359 425581 251397
rect 425481 251325 425497 251359
rect 425565 251325 425581 251359
rect 425481 251309 425581 251325
rect 425757 251359 425857 251397
rect 425757 251325 425773 251359
rect 425841 251325 425857 251359
rect 425757 251309 425857 251325
rect 426033 251359 426133 251397
rect 426033 251325 426049 251359
rect 426117 251325 426133 251359
rect 426033 251309 426133 251325
rect 426309 251359 426409 251397
rect 426309 251325 426325 251359
rect 426393 251325 426409 251359
rect 426309 251309 426409 251325
rect 426585 251359 426685 251397
rect 426585 251325 426601 251359
rect 426669 251325 426685 251359
rect 426585 251309 426685 251325
rect 426861 251359 426961 251397
rect 426861 251325 426877 251359
rect 426945 251325 426961 251359
rect 426861 251309 426961 251325
rect 427137 251359 427237 251397
rect 427137 251325 427153 251359
rect 427221 251325 427237 251359
rect 427137 251309 427237 251325
rect 503337 251553 503437 251569
rect 503337 251519 503353 251553
rect 503421 251519 503437 251553
rect 503337 251481 503437 251519
rect 503613 251553 503713 251569
rect 503613 251519 503629 251553
rect 503697 251519 503713 251553
rect 503613 251481 503713 251519
rect 503889 251553 503989 251569
rect 503889 251519 503905 251553
rect 503973 251519 503989 251553
rect 503889 251481 503989 251519
rect 504165 251553 504265 251569
rect 504165 251519 504181 251553
rect 504249 251519 504265 251553
rect 504165 251481 504265 251519
rect 504441 251553 504541 251569
rect 504441 251519 504457 251553
rect 504525 251519 504541 251553
rect 504441 251481 504541 251519
rect 504717 251553 504817 251569
rect 504717 251519 504733 251553
rect 504801 251519 504817 251553
rect 504717 251481 504817 251519
rect 504993 251553 505093 251569
rect 504993 251519 505009 251553
rect 505077 251519 505093 251553
rect 504993 251481 505093 251519
rect 505269 251553 505369 251569
rect 505269 251519 505285 251553
rect 505353 251519 505369 251553
rect 505269 251481 505369 251519
rect 505545 251553 505645 251569
rect 505545 251519 505561 251553
rect 505629 251519 505645 251553
rect 505545 251481 505645 251519
rect 505821 251553 505921 251569
rect 505821 251519 505837 251553
rect 505905 251519 505921 251553
rect 505821 251481 505921 251519
rect 506097 251553 506197 251569
rect 506097 251519 506113 251553
rect 506181 251519 506197 251553
rect 506097 251481 506197 251519
rect 506373 251553 506473 251569
rect 506373 251519 506389 251553
rect 506457 251519 506473 251553
rect 506373 251481 506473 251519
rect 506649 251553 506749 251569
rect 506649 251519 506665 251553
rect 506733 251519 506749 251553
rect 506649 251481 506749 251519
rect 506925 251553 507025 251569
rect 506925 251519 506941 251553
rect 507009 251519 507025 251553
rect 506925 251481 507025 251519
rect 507201 251553 507301 251569
rect 507201 251519 507217 251553
rect 507285 251519 507301 251553
rect 507201 251481 507301 251519
rect 507477 251553 507577 251569
rect 507477 251519 507493 251553
rect 507561 251519 507577 251553
rect 507477 251481 507577 251519
rect 507753 251553 507853 251569
rect 507753 251519 507769 251553
rect 507837 251519 507853 251553
rect 507753 251481 507853 251519
rect 508029 251553 508129 251569
rect 508029 251519 508045 251553
rect 508113 251519 508129 251553
rect 508029 251481 508129 251519
rect 508305 251553 508405 251569
rect 508305 251519 508321 251553
rect 508389 251519 508405 251553
rect 508305 251481 508405 251519
rect 508581 251553 508681 251569
rect 508581 251519 508597 251553
rect 508665 251519 508681 251553
rect 508581 251481 508681 251519
rect 508857 251553 508957 251569
rect 508857 251519 508873 251553
rect 508941 251519 508957 251553
rect 508857 251481 508957 251519
rect 509133 251553 509233 251569
rect 509133 251519 509149 251553
rect 509217 251519 509233 251553
rect 509133 251481 509233 251519
rect 509409 251553 509509 251569
rect 509409 251519 509425 251553
rect 509493 251519 509509 251553
rect 509409 251481 509509 251519
rect 509685 251553 509785 251569
rect 509685 251519 509701 251553
rect 509769 251519 509785 251553
rect 509685 251481 509785 251519
rect 509961 251553 510061 251569
rect 509961 251519 509977 251553
rect 510045 251519 510061 251553
rect 509961 251481 510061 251519
rect 510237 251553 510337 251569
rect 510237 251519 510253 251553
rect 510321 251519 510337 251553
rect 510237 251481 510337 251519
rect 510513 251553 510613 251569
rect 510513 251519 510529 251553
rect 510597 251519 510613 251553
rect 510513 251481 510613 251519
rect 510789 251553 510889 251569
rect 510789 251519 510805 251553
rect 510873 251519 510889 251553
rect 510789 251481 510889 251519
rect 511065 251553 511165 251569
rect 511065 251519 511081 251553
rect 511149 251519 511165 251553
rect 511065 251481 511165 251519
rect 511341 251553 511441 251569
rect 511341 251519 511357 251553
rect 511425 251519 511441 251553
rect 511341 251481 511441 251519
rect 511617 251553 511717 251569
rect 511617 251519 511633 251553
rect 511701 251519 511717 251553
rect 511617 251481 511717 251519
rect 511893 251553 511993 251569
rect 511893 251519 511909 251553
rect 511977 251519 511993 251553
rect 511893 251481 511993 251519
rect 512169 251553 512269 251569
rect 512169 251519 512185 251553
rect 512253 251519 512269 251553
rect 512169 251481 512269 251519
rect 512445 251553 512545 251569
rect 512445 251519 512461 251553
rect 512529 251519 512545 251553
rect 512445 251481 512545 251519
rect 512721 251553 512821 251569
rect 512721 251519 512737 251553
rect 512805 251519 512821 251553
rect 512721 251481 512821 251519
rect 512997 251553 513097 251569
rect 512997 251519 513013 251553
rect 513081 251519 513097 251553
rect 512997 251481 513097 251519
rect 513273 251553 513373 251569
rect 513273 251519 513289 251553
rect 513357 251519 513373 251553
rect 513273 251481 513373 251519
rect 513549 251553 513649 251569
rect 513549 251519 513565 251553
rect 513633 251519 513649 251553
rect 513549 251481 513649 251519
rect 513825 251553 513925 251569
rect 513825 251519 513841 251553
rect 513909 251519 513925 251553
rect 513825 251481 513925 251519
rect 514101 251553 514201 251569
rect 514101 251519 514117 251553
rect 514185 251519 514201 251553
rect 514101 251481 514201 251519
rect 514377 251553 514477 251569
rect 514377 251519 514393 251553
rect 514461 251519 514477 251553
rect 514377 251481 514477 251519
rect 514653 251553 514753 251569
rect 514653 251519 514669 251553
rect 514737 251519 514753 251553
rect 514653 251481 514753 251519
rect 514929 251553 515029 251569
rect 514929 251519 514945 251553
rect 515013 251519 515029 251553
rect 514929 251481 515029 251519
rect 515205 251553 515305 251569
rect 515205 251519 515221 251553
rect 515289 251519 515305 251553
rect 515205 251481 515305 251519
rect 515481 251553 515581 251569
rect 515481 251519 515497 251553
rect 515565 251519 515581 251553
rect 515481 251481 515581 251519
rect 515757 251553 515857 251569
rect 515757 251519 515773 251553
rect 515841 251519 515857 251553
rect 515757 251481 515857 251519
rect 516033 251553 516133 251569
rect 516033 251519 516049 251553
rect 516117 251519 516133 251553
rect 516033 251481 516133 251519
rect 516309 251553 516409 251569
rect 516309 251519 516325 251553
rect 516393 251519 516409 251553
rect 516309 251481 516409 251519
rect 516585 251553 516685 251569
rect 516585 251519 516601 251553
rect 516669 251519 516685 251553
rect 516585 251481 516685 251519
rect 516861 251553 516961 251569
rect 516861 251519 516877 251553
rect 516945 251519 516961 251553
rect 516861 251481 516961 251519
rect 517137 251553 517237 251569
rect 517137 251519 517153 251553
rect 517221 251519 517237 251553
rect 517137 251481 517237 251519
rect 503337 251359 503437 251397
rect 503337 251325 503353 251359
rect 503421 251325 503437 251359
rect 503337 251309 503437 251325
rect 503613 251359 503713 251397
rect 503613 251325 503629 251359
rect 503697 251325 503713 251359
rect 503613 251309 503713 251325
rect 503889 251359 503989 251397
rect 503889 251325 503905 251359
rect 503973 251325 503989 251359
rect 503889 251309 503989 251325
rect 504165 251359 504265 251397
rect 504165 251325 504181 251359
rect 504249 251325 504265 251359
rect 504165 251309 504265 251325
rect 504441 251359 504541 251397
rect 504441 251325 504457 251359
rect 504525 251325 504541 251359
rect 504441 251309 504541 251325
rect 504717 251359 504817 251397
rect 504717 251325 504733 251359
rect 504801 251325 504817 251359
rect 504717 251309 504817 251325
rect 504993 251359 505093 251397
rect 504993 251325 505009 251359
rect 505077 251325 505093 251359
rect 504993 251309 505093 251325
rect 505269 251359 505369 251397
rect 505269 251325 505285 251359
rect 505353 251325 505369 251359
rect 505269 251309 505369 251325
rect 505545 251359 505645 251397
rect 505545 251325 505561 251359
rect 505629 251325 505645 251359
rect 505545 251309 505645 251325
rect 505821 251359 505921 251397
rect 505821 251325 505837 251359
rect 505905 251325 505921 251359
rect 505821 251309 505921 251325
rect 506097 251359 506197 251397
rect 506097 251325 506113 251359
rect 506181 251325 506197 251359
rect 506097 251309 506197 251325
rect 506373 251359 506473 251397
rect 506373 251325 506389 251359
rect 506457 251325 506473 251359
rect 506373 251309 506473 251325
rect 506649 251359 506749 251397
rect 506649 251325 506665 251359
rect 506733 251325 506749 251359
rect 506649 251309 506749 251325
rect 506925 251359 507025 251397
rect 506925 251325 506941 251359
rect 507009 251325 507025 251359
rect 506925 251309 507025 251325
rect 507201 251359 507301 251397
rect 507201 251325 507217 251359
rect 507285 251325 507301 251359
rect 507201 251309 507301 251325
rect 507477 251359 507577 251397
rect 507477 251325 507493 251359
rect 507561 251325 507577 251359
rect 507477 251309 507577 251325
rect 507753 251359 507853 251397
rect 507753 251325 507769 251359
rect 507837 251325 507853 251359
rect 507753 251309 507853 251325
rect 508029 251359 508129 251397
rect 508029 251325 508045 251359
rect 508113 251325 508129 251359
rect 508029 251309 508129 251325
rect 508305 251359 508405 251397
rect 508305 251325 508321 251359
rect 508389 251325 508405 251359
rect 508305 251309 508405 251325
rect 508581 251359 508681 251397
rect 508581 251325 508597 251359
rect 508665 251325 508681 251359
rect 508581 251309 508681 251325
rect 508857 251359 508957 251397
rect 508857 251325 508873 251359
rect 508941 251325 508957 251359
rect 508857 251309 508957 251325
rect 509133 251359 509233 251397
rect 509133 251325 509149 251359
rect 509217 251325 509233 251359
rect 509133 251309 509233 251325
rect 509409 251359 509509 251397
rect 509409 251325 509425 251359
rect 509493 251325 509509 251359
rect 509409 251309 509509 251325
rect 509685 251359 509785 251397
rect 509685 251325 509701 251359
rect 509769 251325 509785 251359
rect 509685 251309 509785 251325
rect 509961 251359 510061 251397
rect 509961 251325 509977 251359
rect 510045 251325 510061 251359
rect 509961 251309 510061 251325
rect 510237 251359 510337 251397
rect 510237 251325 510253 251359
rect 510321 251325 510337 251359
rect 510237 251309 510337 251325
rect 510513 251359 510613 251397
rect 510513 251325 510529 251359
rect 510597 251325 510613 251359
rect 510513 251309 510613 251325
rect 510789 251359 510889 251397
rect 510789 251325 510805 251359
rect 510873 251325 510889 251359
rect 510789 251309 510889 251325
rect 511065 251359 511165 251397
rect 511065 251325 511081 251359
rect 511149 251325 511165 251359
rect 511065 251309 511165 251325
rect 511341 251359 511441 251397
rect 511341 251325 511357 251359
rect 511425 251325 511441 251359
rect 511341 251309 511441 251325
rect 511617 251359 511717 251397
rect 511617 251325 511633 251359
rect 511701 251325 511717 251359
rect 511617 251309 511717 251325
rect 511893 251359 511993 251397
rect 511893 251325 511909 251359
rect 511977 251325 511993 251359
rect 511893 251309 511993 251325
rect 512169 251359 512269 251397
rect 512169 251325 512185 251359
rect 512253 251325 512269 251359
rect 512169 251309 512269 251325
rect 512445 251359 512545 251397
rect 512445 251325 512461 251359
rect 512529 251325 512545 251359
rect 512445 251309 512545 251325
rect 512721 251359 512821 251397
rect 512721 251325 512737 251359
rect 512805 251325 512821 251359
rect 512721 251309 512821 251325
rect 512997 251359 513097 251397
rect 512997 251325 513013 251359
rect 513081 251325 513097 251359
rect 512997 251309 513097 251325
rect 513273 251359 513373 251397
rect 513273 251325 513289 251359
rect 513357 251325 513373 251359
rect 513273 251309 513373 251325
rect 513549 251359 513649 251397
rect 513549 251325 513565 251359
rect 513633 251325 513649 251359
rect 513549 251309 513649 251325
rect 513825 251359 513925 251397
rect 513825 251325 513841 251359
rect 513909 251325 513925 251359
rect 513825 251309 513925 251325
rect 514101 251359 514201 251397
rect 514101 251325 514117 251359
rect 514185 251325 514201 251359
rect 514101 251309 514201 251325
rect 514377 251359 514477 251397
rect 514377 251325 514393 251359
rect 514461 251325 514477 251359
rect 514377 251309 514477 251325
rect 514653 251359 514753 251397
rect 514653 251325 514669 251359
rect 514737 251325 514753 251359
rect 514653 251309 514753 251325
rect 514929 251359 515029 251397
rect 514929 251325 514945 251359
rect 515013 251325 515029 251359
rect 514929 251309 515029 251325
rect 515205 251359 515305 251397
rect 515205 251325 515221 251359
rect 515289 251325 515305 251359
rect 515205 251309 515305 251325
rect 515481 251359 515581 251397
rect 515481 251325 515497 251359
rect 515565 251325 515581 251359
rect 515481 251309 515581 251325
rect 515757 251359 515857 251397
rect 515757 251325 515773 251359
rect 515841 251325 515857 251359
rect 515757 251309 515857 251325
rect 516033 251359 516133 251397
rect 516033 251325 516049 251359
rect 516117 251325 516133 251359
rect 516033 251309 516133 251325
rect 516309 251359 516409 251397
rect 516309 251325 516325 251359
rect 516393 251325 516409 251359
rect 516309 251309 516409 251325
rect 516585 251359 516685 251397
rect 516585 251325 516601 251359
rect 516669 251325 516685 251359
rect 516585 251309 516685 251325
rect 516861 251359 516961 251397
rect 516861 251325 516877 251359
rect 516945 251325 516961 251359
rect 516861 251309 516961 251325
rect 517137 251359 517237 251397
rect 517137 251325 517153 251359
rect 517221 251325 517237 251359
rect 517137 251309 517237 251325
rect 322694 250957 322794 250973
rect 322694 250923 322710 250957
rect 322778 250923 322794 250957
rect 322694 250885 322794 250923
rect 322970 250957 323070 250973
rect 322970 250923 322986 250957
rect 323054 250923 323070 250957
rect 322970 250885 323070 250923
rect 323246 250957 323346 250973
rect 323246 250923 323262 250957
rect 323330 250923 323346 250957
rect 323246 250885 323346 250923
rect 323522 250957 323622 250973
rect 323522 250923 323538 250957
rect 323606 250923 323622 250957
rect 323522 250885 323622 250923
rect 323798 250957 323898 250973
rect 323798 250923 323814 250957
rect 323882 250923 323898 250957
rect 323798 250885 323898 250923
rect 324074 250957 324174 250973
rect 324074 250923 324090 250957
rect 324158 250923 324174 250957
rect 324074 250885 324174 250923
rect 324350 250957 324450 250973
rect 324350 250923 324366 250957
rect 324434 250923 324450 250957
rect 324350 250885 324450 250923
rect 324626 250957 324726 250973
rect 324626 250923 324642 250957
rect 324710 250923 324726 250957
rect 324626 250885 324726 250923
rect 324902 250957 325002 250973
rect 324902 250923 324918 250957
rect 324986 250923 325002 250957
rect 324902 250885 325002 250923
rect 325178 250957 325278 250973
rect 325178 250923 325194 250957
rect 325262 250923 325278 250957
rect 325178 250885 325278 250923
rect 325454 250957 325554 250973
rect 325454 250923 325470 250957
rect 325538 250923 325554 250957
rect 325454 250885 325554 250923
rect 325730 250957 325830 250973
rect 325730 250923 325746 250957
rect 325814 250923 325830 250957
rect 325730 250885 325830 250923
rect 326006 250957 326106 250973
rect 326006 250923 326022 250957
rect 326090 250923 326106 250957
rect 326006 250885 326106 250923
rect 326282 250957 326382 250973
rect 326282 250923 326298 250957
rect 326366 250923 326382 250957
rect 326282 250885 326382 250923
rect 326558 250957 326658 250973
rect 326558 250923 326574 250957
rect 326642 250923 326658 250957
rect 326558 250885 326658 250923
rect 326834 250957 326934 250973
rect 326834 250923 326850 250957
rect 326918 250923 326934 250957
rect 326834 250885 326934 250923
rect 327110 250957 327210 250973
rect 327110 250923 327126 250957
rect 327194 250923 327210 250957
rect 327110 250885 327210 250923
rect 327386 250957 327486 250973
rect 327386 250923 327402 250957
rect 327470 250923 327486 250957
rect 327386 250885 327486 250923
rect 327662 250957 327762 250973
rect 327662 250923 327678 250957
rect 327746 250923 327762 250957
rect 327662 250885 327762 250923
rect 327938 250957 328038 250973
rect 327938 250923 327954 250957
rect 328022 250923 328038 250957
rect 327938 250885 328038 250923
rect 328214 250957 328314 250973
rect 328214 250923 328230 250957
rect 328298 250923 328314 250957
rect 328214 250885 328314 250923
rect 328490 250957 328590 250973
rect 328490 250923 328506 250957
rect 328574 250923 328590 250957
rect 328490 250885 328590 250923
rect 328766 250957 328866 250973
rect 328766 250923 328782 250957
rect 328850 250923 328866 250957
rect 328766 250885 328866 250923
rect 329042 250957 329142 250973
rect 329042 250923 329058 250957
rect 329126 250923 329142 250957
rect 329042 250885 329142 250923
rect 329318 250957 329418 250973
rect 329318 250923 329334 250957
rect 329402 250923 329418 250957
rect 329318 250885 329418 250923
rect 329594 250957 329694 250973
rect 329594 250923 329610 250957
rect 329678 250923 329694 250957
rect 329594 250885 329694 250923
rect 329870 250957 329970 250973
rect 329870 250923 329886 250957
rect 329954 250923 329970 250957
rect 329870 250885 329970 250923
rect 330146 250957 330246 250973
rect 330146 250923 330162 250957
rect 330230 250923 330246 250957
rect 330146 250885 330246 250923
rect 330422 250957 330522 250973
rect 330422 250923 330438 250957
rect 330506 250923 330522 250957
rect 330422 250885 330522 250923
rect 330698 250957 330798 250973
rect 330698 250923 330714 250957
rect 330782 250923 330798 250957
rect 330698 250885 330798 250923
rect 330974 250957 331074 250973
rect 330974 250923 330990 250957
rect 331058 250923 331074 250957
rect 330974 250885 331074 250923
rect 331250 250957 331350 250973
rect 331250 250923 331266 250957
rect 331334 250923 331350 250957
rect 331250 250885 331350 250923
rect 331526 250957 331626 250973
rect 331526 250923 331542 250957
rect 331610 250923 331626 250957
rect 331526 250885 331626 250923
rect 331802 250957 331902 250973
rect 331802 250923 331818 250957
rect 331886 250923 331902 250957
rect 331802 250885 331902 250923
rect 332078 250957 332178 250973
rect 332078 250923 332094 250957
rect 332162 250923 332178 250957
rect 332078 250885 332178 250923
rect 332354 250957 332454 250973
rect 332354 250923 332370 250957
rect 332438 250923 332454 250957
rect 332354 250885 332454 250923
rect 332630 250957 332730 250973
rect 332630 250923 332646 250957
rect 332714 250923 332730 250957
rect 332630 250885 332730 250923
rect 332906 250957 333006 250973
rect 332906 250923 332922 250957
rect 332990 250923 333006 250957
rect 332906 250885 333006 250923
rect 333182 250957 333282 250973
rect 333182 250923 333198 250957
rect 333266 250923 333282 250957
rect 333182 250885 333282 250923
rect 333458 250957 333558 250973
rect 333458 250923 333474 250957
rect 333542 250923 333558 250957
rect 333458 250885 333558 250923
rect 333734 250957 333834 250973
rect 333734 250923 333750 250957
rect 333818 250923 333834 250957
rect 333734 250885 333834 250923
rect 334010 250957 334110 250973
rect 334010 250923 334026 250957
rect 334094 250923 334110 250957
rect 334010 250885 334110 250923
rect 334286 250957 334386 250973
rect 334286 250923 334302 250957
rect 334370 250923 334386 250957
rect 334286 250885 334386 250923
rect 334562 250957 334662 250973
rect 334562 250923 334578 250957
rect 334646 250923 334662 250957
rect 334562 250885 334662 250923
rect 334838 250957 334938 250973
rect 334838 250923 334854 250957
rect 334922 250923 334938 250957
rect 334838 250885 334938 250923
rect 335114 250957 335214 250973
rect 335114 250923 335130 250957
rect 335198 250923 335214 250957
rect 335114 250885 335214 250923
rect 335390 250957 335490 250973
rect 335390 250923 335406 250957
rect 335474 250923 335490 250957
rect 335390 250885 335490 250923
rect 335666 250957 335766 250973
rect 335666 250923 335682 250957
rect 335750 250923 335766 250957
rect 335666 250885 335766 250923
rect 335942 250957 336042 250973
rect 335942 250923 335958 250957
rect 336026 250923 336042 250957
rect 335942 250885 336042 250923
rect 336218 250957 336318 250973
rect 336218 250923 336234 250957
rect 336302 250923 336318 250957
rect 336218 250885 336318 250923
rect 336494 250957 336594 250973
rect 336494 250923 336510 250957
rect 336578 250923 336594 250957
rect 336494 250885 336594 250923
rect 322694 250763 322794 250801
rect 322694 250729 322710 250763
rect 322778 250729 322794 250763
rect 322694 250713 322794 250729
rect 322970 250763 323070 250801
rect 322970 250729 322986 250763
rect 323054 250729 323070 250763
rect 322970 250713 323070 250729
rect 323246 250763 323346 250801
rect 323246 250729 323262 250763
rect 323330 250729 323346 250763
rect 323246 250713 323346 250729
rect 323522 250763 323622 250801
rect 323522 250729 323538 250763
rect 323606 250729 323622 250763
rect 323522 250713 323622 250729
rect 323798 250763 323898 250801
rect 323798 250729 323814 250763
rect 323882 250729 323898 250763
rect 323798 250713 323898 250729
rect 324074 250763 324174 250801
rect 324074 250729 324090 250763
rect 324158 250729 324174 250763
rect 324074 250713 324174 250729
rect 324350 250763 324450 250801
rect 324350 250729 324366 250763
rect 324434 250729 324450 250763
rect 324350 250713 324450 250729
rect 324626 250763 324726 250801
rect 324626 250729 324642 250763
rect 324710 250729 324726 250763
rect 324626 250713 324726 250729
rect 324902 250763 325002 250801
rect 324902 250729 324918 250763
rect 324986 250729 325002 250763
rect 324902 250713 325002 250729
rect 325178 250763 325278 250801
rect 325178 250729 325194 250763
rect 325262 250729 325278 250763
rect 325178 250713 325278 250729
rect 325454 250763 325554 250801
rect 325454 250729 325470 250763
rect 325538 250729 325554 250763
rect 325454 250713 325554 250729
rect 325730 250763 325830 250801
rect 325730 250729 325746 250763
rect 325814 250729 325830 250763
rect 325730 250713 325830 250729
rect 326006 250763 326106 250801
rect 326006 250729 326022 250763
rect 326090 250729 326106 250763
rect 326006 250713 326106 250729
rect 326282 250763 326382 250801
rect 326282 250729 326298 250763
rect 326366 250729 326382 250763
rect 326282 250713 326382 250729
rect 326558 250763 326658 250801
rect 326558 250729 326574 250763
rect 326642 250729 326658 250763
rect 326558 250713 326658 250729
rect 326834 250763 326934 250801
rect 326834 250729 326850 250763
rect 326918 250729 326934 250763
rect 326834 250713 326934 250729
rect 327110 250763 327210 250801
rect 327110 250729 327126 250763
rect 327194 250729 327210 250763
rect 327110 250713 327210 250729
rect 327386 250763 327486 250801
rect 327386 250729 327402 250763
rect 327470 250729 327486 250763
rect 327386 250713 327486 250729
rect 327662 250763 327762 250801
rect 327662 250729 327678 250763
rect 327746 250729 327762 250763
rect 327662 250713 327762 250729
rect 327938 250763 328038 250801
rect 327938 250729 327954 250763
rect 328022 250729 328038 250763
rect 327938 250713 328038 250729
rect 328214 250763 328314 250801
rect 328214 250729 328230 250763
rect 328298 250729 328314 250763
rect 328214 250713 328314 250729
rect 328490 250763 328590 250801
rect 328490 250729 328506 250763
rect 328574 250729 328590 250763
rect 328490 250713 328590 250729
rect 328766 250763 328866 250801
rect 328766 250729 328782 250763
rect 328850 250729 328866 250763
rect 328766 250713 328866 250729
rect 329042 250763 329142 250801
rect 329042 250729 329058 250763
rect 329126 250729 329142 250763
rect 329042 250713 329142 250729
rect 329318 250763 329418 250801
rect 329318 250729 329334 250763
rect 329402 250729 329418 250763
rect 329318 250713 329418 250729
rect 329594 250763 329694 250801
rect 329594 250729 329610 250763
rect 329678 250729 329694 250763
rect 329594 250713 329694 250729
rect 329870 250763 329970 250801
rect 329870 250729 329886 250763
rect 329954 250729 329970 250763
rect 329870 250713 329970 250729
rect 330146 250763 330246 250801
rect 330146 250729 330162 250763
rect 330230 250729 330246 250763
rect 330146 250713 330246 250729
rect 330422 250763 330522 250801
rect 330422 250729 330438 250763
rect 330506 250729 330522 250763
rect 330422 250713 330522 250729
rect 330698 250763 330798 250801
rect 330698 250729 330714 250763
rect 330782 250729 330798 250763
rect 330698 250713 330798 250729
rect 330974 250763 331074 250801
rect 330974 250729 330990 250763
rect 331058 250729 331074 250763
rect 330974 250713 331074 250729
rect 331250 250763 331350 250801
rect 331250 250729 331266 250763
rect 331334 250729 331350 250763
rect 331250 250713 331350 250729
rect 331526 250763 331626 250801
rect 331526 250729 331542 250763
rect 331610 250729 331626 250763
rect 331526 250713 331626 250729
rect 331802 250763 331902 250801
rect 331802 250729 331818 250763
rect 331886 250729 331902 250763
rect 331802 250713 331902 250729
rect 332078 250763 332178 250801
rect 332078 250729 332094 250763
rect 332162 250729 332178 250763
rect 332078 250713 332178 250729
rect 332354 250763 332454 250801
rect 332354 250729 332370 250763
rect 332438 250729 332454 250763
rect 332354 250713 332454 250729
rect 332630 250763 332730 250801
rect 332630 250729 332646 250763
rect 332714 250729 332730 250763
rect 332630 250713 332730 250729
rect 332906 250763 333006 250801
rect 332906 250729 332922 250763
rect 332990 250729 333006 250763
rect 332906 250713 333006 250729
rect 333182 250763 333282 250801
rect 333182 250729 333198 250763
rect 333266 250729 333282 250763
rect 333182 250713 333282 250729
rect 333458 250763 333558 250801
rect 333458 250729 333474 250763
rect 333542 250729 333558 250763
rect 333458 250713 333558 250729
rect 333734 250763 333834 250801
rect 333734 250729 333750 250763
rect 333818 250729 333834 250763
rect 333734 250713 333834 250729
rect 334010 250763 334110 250801
rect 334010 250729 334026 250763
rect 334094 250729 334110 250763
rect 334010 250713 334110 250729
rect 334286 250763 334386 250801
rect 334286 250729 334302 250763
rect 334370 250729 334386 250763
rect 334286 250713 334386 250729
rect 334562 250763 334662 250801
rect 334562 250729 334578 250763
rect 334646 250729 334662 250763
rect 334562 250713 334662 250729
rect 334838 250763 334938 250801
rect 334838 250729 334854 250763
rect 334922 250729 334938 250763
rect 334838 250713 334938 250729
rect 335114 250763 335214 250801
rect 335114 250729 335130 250763
rect 335198 250729 335214 250763
rect 335114 250713 335214 250729
rect 335390 250763 335490 250801
rect 335390 250729 335406 250763
rect 335474 250729 335490 250763
rect 335390 250713 335490 250729
rect 335666 250763 335766 250801
rect 335666 250729 335682 250763
rect 335750 250729 335766 250763
rect 335666 250713 335766 250729
rect 335942 250763 336042 250801
rect 335942 250729 335958 250763
rect 336026 250729 336042 250763
rect 335942 250713 336042 250729
rect 336218 250763 336318 250801
rect 336218 250729 336234 250763
rect 336302 250729 336318 250763
rect 336218 250713 336318 250729
rect 336494 250763 336594 250801
rect 336494 250729 336510 250763
rect 336578 250729 336594 250763
rect 336494 250713 336594 250729
rect 59323 146027 59389 146043
rect 59323 145993 59339 146027
rect 59373 145993 59389 146027
rect 59323 145977 59389 145993
rect 59341 145946 59371 145977
rect 59341 145715 59371 145746
rect 59323 145699 59389 145715
rect 59323 145665 59339 145699
rect 59373 145665 59389 145699
rect 59323 145649 59389 145665
rect 149521 145623 149621 145639
rect 149521 145589 149537 145623
rect 149605 145589 149621 145623
rect 149521 145542 149621 145589
rect 149521 145295 149621 145342
rect 149521 145261 149537 145295
rect 149605 145261 149621 145295
rect 149521 145245 149621 145261
rect 239340 146056 239406 146072
rect 239340 146022 239356 146056
rect 239390 146022 239406 146056
rect 239340 146006 239406 146022
rect 239358 145984 239388 146006
rect 239358 145762 239388 145784
rect 239340 145746 239406 145762
rect 239340 145712 239356 145746
rect 239390 145712 239406 145746
rect 239340 145696 239406 145712
rect 329323 146027 329389 146043
rect 329323 145993 329339 146027
rect 329373 145993 329389 146027
rect 329323 145977 329389 145993
rect 329341 145946 329371 145977
rect 329341 145715 329371 145746
rect 329323 145699 329389 145715
rect 329323 145665 329339 145699
rect 329373 145665 329389 145699
rect 329323 145649 329389 145665
rect 419521 145623 419621 145639
rect 419521 145589 419537 145623
rect 419605 145589 419621 145623
rect 419521 145542 419621 145589
rect 419521 145295 419621 145342
rect 419521 145261 419537 145295
rect 419605 145261 419621 145295
rect 419521 145245 419621 145261
rect 509340 146056 509406 146072
rect 509340 146022 509356 146056
rect 509390 146022 509406 146056
rect 509340 146006 509406 146022
rect 509358 145984 509388 146006
rect 509358 145762 509388 145784
rect 509340 145746 509406 145762
rect 509340 145712 509356 145746
rect 509390 145712 509406 145746
rect 509340 145696 509406 145712
rect 59340 56056 59406 56072
rect 59340 56022 59356 56056
rect 59390 56022 59406 56056
rect 59340 56006 59406 56022
rect 59358 55984 59388 56006
rect 59358 55762 59388 55784
rect 59340 55746 59406 55762
rect 59340 55712 59356 55746
rect 59390 55712 59406 55746
rect 59340 55696 59406 55712
rect 149611 56055 149711 56071
rect 149611 56021 149627 56055
rect 149695 56021 149711 56055
rect 149611 55983 149711 56021
rect 149611 55745 149711 55783
rect 149611 55711 149627 55745
rect 149695 55711 149711 55745
rect 149611 55695 149711 55711
rect 239621 55765 239721 55781
rect 239621 55731 239637 55765
rect 239705 55731 239721 55765
rect 239621 55693 239721 55731
rect 239621 55455 239721 55493
rect 239621 55421 239637 55455
rect 239705 55421 239721 55455
rect 239621 55405 239721 55421
rect 329340 56056 329406 56072
rect 329340 56022 329356 56056
rect 329390 56022 329406 56056
rect 329340 56006 329406 56022
rect 329358 55984 329388 56006
rect 329358 55762 329388 55784
rect 329340 55746 329406 55762
rect 329340 55712 329356 55746
rect 329390 55712 329406 55746
rect 329340 55696 329406 55712
rect 419611 56055 419711 56071
rect 419611 56021 419627 56055
rect 419695 56021 419711 56055
rect 419611 55983 419711 56021
rect 419611 55745 419711 55783
rect 419611 55711 419627 55745
rect 419695 55711 419711 55745
rect 419611 55695 419711 55711
rect 509621 55765 509721 55781
rect 509621 55731 509637 55765
rect 509705 55731 509721 55765
rect 509621 55693 509721 55731
rect 509621 55455 509721 55493
rect 509621 55421 509637 55455
rect 509705 55421 509721 55455
rect 509621 55405 509721 55421
<< polycont >>
rect 329158 657946 329192 657980
rect 329158 657636 329192 657670
rect 419339 657513 419407 657547
rect 419339 657185 419407 657219
rect 509158 657946 509192 657980
rect 509158 657636 509192 657670
rect 59627 656021 59695 656055
rect 59627 655711 59695 655745
rect 149356 656022 149390 656056
rect 149356 655712 149390 655746
rect 239339 655993 239373 656027
rect 239339 655665 239373 655699
rect 419429 582945 419497 582979
rect 419429 582635 419497 582669
rect 509439 582655 509507 582689
rect 509439 582345 509507 582379
rect 59627 581021 59695 581055
rect 59627 580711 59695 580745
rect 149637 580731 149705 580765
rect 149637 580421 149705 580455
rect 239356 581022 239390 581056
rect 239356 580712 239390 580746
rect 329537 580589 329605 580623
rect 329537 580261 329605 580295
rect 58903 491809 58971 491843
rect 59179 491809 59247 491843
rect 59455 491809 59523 491843
rect 59731 491809 59799 491843
rect 60007 491809 60075 491843
rect 60283 491809 60351 491843
rect 60559 491809 60627 491843
rect 60835 491809 60903 491843
rect 61111 491809 61179 491843
rect 61387 491809 61455 491843
rect 58903 491615 58971 491649
rect 59179 491615 59247 491649
rect 59455 491615 59523 491649
rect 59731 491615 59799 491649
rect 60007 491615 60075 491649
rect 60283 491615 60351 491649
rect 60559 491615 60627 491649
rect 60835 491615 60903 491649
rect 61111 491615 61179 491649
rect 61387 491615 61455 491649
rect 323893 492197 323961 492231
rect 324169 492197 324237 492231
rect 324445 492197 324513 492231
rect 324721 492197 324789 492231
rect 324997 492197 325065 492231
rect 325273 492197 325341 492231
rect 325549 492197 325617 492231
rect 325825 492197 325893 492231
rect 326101 492197 326169 492231
rect 326377 492197 326445 492231
rect 326653 492197 326721 492231
rect 326929 492197 326997 492231
rect 327205 492197 327273 492231
rect 327481 492197 327549 492231
rect 327757 492197 327825 492231
rect 328033 492197 328101 492231
rect 328309 492197 328377 492231
rect 328585 492197 328653 492231
rect 328861 492197 328929 492231
rect 329137 492197 329205 492231
rect 329413 492197 329481 492231
rect 329689 492197 329757 492231
rect 329965 492197 330033 492231
rect 330241 492197 330309 492231
rect 330517 492197 330585 492231
rect 330793 492197 330861 492231
rect 331069 492197 331137 492231
rect 331345 492197 331413 492231
rect 331621 492197 331689 492231
rect 331897 492197 331965 492231
rect 332173 492197 332241 492231
rect 332449 492197 332517 492231
rect 332725 492197 332793 492231
rect 333001 492197 333069 492231
rect 333277 492197 333345 492231
rect 333553 492197 333621 492231
rect 333829 492197 333897 492231
rect 334105 492197 334173 492231
rect 334381 492197 334449 492231
rect 334657 492197 334725 492231
rect 334933 492197 335001 492231
rect 335209 492197 335277 492231
rect 335485 492197 335553 492231
rect 335761 492197 335829 492231
rect 336037 492197 336105 492231
rect 336313 492197 336381 492231
rect 336589 492197 336657 492231
rect 336865 492197 336933 492231
rect 337141 492197 337209 492231
rect 337417 492197 337485 492231
rect 337693 492197 337761 492231
rect 323893 492003 323961 492037
rect 324169 492003 324237 492037
rect 324445 492003 324513 492037
rect 324721 492003 324789 492037
rect 324997 492003 325065 492037
rect 325273 492003 325341 492037
rect 325549 492003 325617 492037
rect 325825 492003 325893 492037
rect 326101 492003 326169 492037
rect 326377 492003 326445 492037
rect 326653 492003 326721 492037
rect 326929 492003 326997 492037
rect 327205 492003 327273 492037
rect 327481 492003 327549 492037
rect 327757 492003 327825 492037
rect 328033 492003 328101 492037
rect 328309 492003 328377 492037
rect 328585 492003 328653 492037
rect 328861 492003 328929 492037
rect 329137 492003 329205 492037
rect 329413 492003 329481 492037
rect 329689 492003 329757 492037
rect 329965 492003 330033 492037
rect 330241 492003 330309 492037
rect 330517 492003 330585 492037
rect 330793 492003 330861 492037
rect 331069 492003 331137 492037
rect 331345 492003 331413 492037
rect 331621 492003 331689 492037
rect 331897 492003 331965 492037
rect 332173 492003 332241 492037
rect 332449 492003 332517 492037
rect 332725 492003 332793 492037
rect 333001 492003 333069 492037
rect 333277 492003 333345 492037
rect 333553 492003 333621 492037
rect 333829 492003 333897 492037
rect 334105 492003 334173 492037
rect 334381 492003 334449 492037
rect 334657 492003 334725 492037
rect 334933 492003 335001 492037
rect 335209 492003 335277 492037
rect 335485 492003 335553 492037
rect 335761 492003 335829 492037
rect 336037 492003 336105 492037
rect 336313 492003 336381 492037
rect 336589 492003 336657 492037
rect 336865 492003 336933 492037
rect 337141 492003 337209 492037
rect 337417 492003 337485 492037
rect 337693 492003 337761 492037
rect 143353 491519 143421 491553
rect 143629 491519 143697 491553
rect 143905 491519 143973 491553
rect 144181 491519 144249 491553
rect 144457 491519 144525 491553
rect 144733 491519 144801 491553
rect 145009 491519 145077 491553
rect 145285 491519 145353 491553
rect 145561 491519 145629 491553
rect 145837 491519 145905 491553
rect 146113 491519 146181 491553
rect 146389 491519 146457 491553
rect 146665 491519 146733 491553
rect 146941 491519 147009 491553
rect 147217 491519 147285 491553
rect 147493 491519 147561 491553
rect 147769 491519 147837 491553
rect 148045 491519 148113 491553
rect 148321 491519 148389 491553
rect 148597 491519 148665 491553
rect 148873 491519 148941 491553
rect 149149 491519 149217 491553
rect 149425 491519 149493 491553
rect 149701 491519 149769 491553
rect 149977 491519 150045 491553
rect 150253 491519 150321 491553
rect 150529 491519 150597 491553
rect 150805 491519 150873 491553
rect 151081 491519 151149 491553
rect 151357 491519 151425 491553
rect 151633 491519 151701 491553
rect 151909 491519 151977 491553
rect 152185 491519 152253 491553
rect 152461 491519 152529 491553
rect 152737 491519 152805 491553
rect 153013 491519 153081 491553
rect 153289 491519 153357 491553
rect 153565 491519 153633 491553
rect 153841 491519 153909 491553
rect 154117 491519 154185 491553
rect 154393 491519 154461 491553
rect 154669 491519 154737 491553
rect 154945 491519 155013 491553
rect 155221 491519 155289 491553
rect 155497 491519 155565 491553
rect 155773 491519 155841 491553
rect 156049 491519 156117 491553
rect 156325 491519 156393 491553
rect 156601 491519 156669 491553
rect 156877 491519 156945 491553
rect 157153 491519 157221 491553
rect 143353 491325 143421 491359
rect 143629 491325 143697 491359
rect 143905 491325 143973 491359
rect 144181 491325 144249 491359
rect 144457 491325 144525 491359
rect 144733 491325 144801 491359
rect 145009 491325 145077 491359
rect 145285 491325 145353 491359
rect 145561 491325 145629 491359
rect 145837 491325 145905 491359
rect 146113 491325 146181 491359
rect 146389 491325 146457 491359
rect 146665 491325 146733 491359
rect 146941 491325 147009 491359
rect 147217 491325 147285 491359
rect 147493 491325 147561 491359
rect 147769 491325 147837 491359
rect 148045 491325 148113 491359
rect 148321 491325 148389 491359
rect 148597 491325 148665 491359
rect 148873 491325 148941 491359
rect 149149 491325 149217 491359
rect 149425 491325 149493 491359
rect 149701 491325 149769 491359
rect 149977 491325 150045 491359
rect 150253 491325 150321 491359
rect 150529 491325 150597 491359
rect 150805 491325 150873 491359
rect 151081 491325 151149 491359
rect 151357 491325 151425 491359
rect 151633 491325 151701 491359
rect 151909 491325 151977 491359
rect 152185 491325 152253 491359
rect 152461 491325 152529 491359
rect 152737 491325 152805 491359
rect 153013 491325 153081 491359
rect 153289 491325 153357 491359
rect 153565 491325 153633 491359
rect 153841 491325 153909 491359
rect 154117 491325 154185 491359
rect 154393 491325 154461 491359
rect 154669 491325 154737 491359
rect 154945 491325 155013 491359
rect 155221 491325 155289 491359
rect 155497 491325 155565 491359
rect 155773 491325 155841 491359
rect 156049 491325 156117 491359
rect 156325 491325 156393 491359
rect 156601 491325 156669 491359
rect 156877 491325 156945 491359
rect 157153 491325 157221 491359
rect 418902 491481 418970 491515
rect 419178 491481 419246 491515
rect 419454 491481 419522 491515
rect 419730 491481 419798 491515
rect 420006 491481 420074 491515
rect 418902 491287 418970 491321
rect 419178 491287 419246 491321
rect 419454 491287 419522 491321
rect 419730 491287 419798 491321
rect 420006 491287 420074 491321
rect 508903 491809 508971 491843
rect 509179 491809 509247 491843
rect 509455 491809 509523 491843
rect 509731 491809 509799 491843
rect 510007 491809 510075 491843
rect 510283 491809 510351 491843
rect 510559 491809 510627 491843
rect 510835 491809 510903 491843
rect 511111 491809 511179 491843
rect 511387 491809 511455 491843
rect 508903 491615 508971 491649
rect 509179 491615 509247 491649
rect 509455 491615 509523 491649
rect 509731 491615 509799 491649
rect 510007 491615 510075 491649
rect 510283 491615 510351 491649
rect 510559 491615 510627 491649
rect 510835 491615 510903 491649
rect 511111 491615 511179 491649
rect 511387 491615 511455 491649
rect 232710 490923 232778 490957
rect 232986 490923 233054 490957
rect 233262 490923 233330 490957
rect 233538 490923 233606 490957
rect 233814 490923 233882 490957
rect 234090 490923 234158 490957
rect 234366 490923 234434 490957
rect 234642 490923 234710 490957
rect 234918 490923 234986 490957
rect 235194 490923 235262 490957
rect 235470 490923 235538 490957
rect 235746 490923 235814 490957
rect 236022 490923 236090 490957
rect 236298 490923 236366 490957
rect 236574 490923 236642 490957
rect 236850 490923 236918 490957
rect 237126 490923 237194 490957
rect 237402 490923 237470 490957
rect 237678 490923 237746 490957
rect 237954 490923 238022 490957
rect 238230 490923 238298 490957
rect 238506 490923 238574 490957
rect 238782 490923 238850 490957
rect 239058 490923 239126 490957
rect 239334 490923 239402 490957
rect 239610 490923 239678 490957
rect 239886 490923 239954 490957
rect 240162 490923 240230 490957
rect 240438 490923 240506 490957
rect 240714 490923 240782 490957
rect 240990 490923 241058 490957
rect 241266 490923 241334 490957
rect 241542 490923 241610 490957
rect 241818 490923 241886 490957
rect 242094 490923 242162 490957
rect 242370 490923 242438 490957
rect 242646 490923 242714 490957
rect 242922 490923 242990 490957
rect 243198 490923 243266 490957
rect 243474 490923 243542 490957
rect 243750 490923 243818 490957
rect 244026 490923 244094 490957
rect 244302 490923 244370 490957
rect 244578 490923 244646 490957
rect 244854 490923 244922 490957
rect 245130 490923 245198 490957
rect 245406 490923 245474 490957
rect 245682 490923 245750 490957
rect 245958 490923 246026 490957
rect 246234 490923 246302 490957
rect 246510 490923 246578 490957
rect 232710 490729 232778 490763
rect 232986 490729 233054 490763
rect 233262 490729 233330 490763
rect 233538 490729 233606 490763
rect 233814 490729 233882 490763
rect 234090 490729 234158 490763
rect 234366 490729 234434 490763
rect 234642 490729 234710 490763
rect 234918 490729 234986 490763
rect 235194 490729 235262 490763
rect 235470 490729 235538 490763
rect 235746 490729 235814 490763
rect 236022 490729 236090 490763
rect 236298 490729 236366 490763
rect 236574 490729 236642 490763
rect 236850 490729 236918 490763
rect 237126 490729 237194 490763
rect 237402 490729 237470 490763
rect 237678 490729 237746 490763
rect 237954 490729 238022 490763
rect 238230 490729 238298 490763
rect 238506 490729 238574 490763
rect 238782 490729 238850 490763
rect 239058 490729 239126 490763
rect 239334 490729 239402 490763
rect 239610 490729 239678 490763
rect 239886 490729 239954 490763
rect 240162 490729 240230 490763
rect 240438 490729 240506 490763
rect 240714 490729 240782 490763
rect 240990 490729 241058 490763
rect 241266 490729 241334 490763
rect 241542 490729 241610 490763
rect 241818 490729 241886 490763
rect 242094 490729 242162 490763
rect 242370 490729 242438 490763
rect 242646 490729 242714 490763
rect 242922 490729 242990 490763
rect 243198 490729 243266 490763
rect 243474 490729 243542 490763
rect 243750 490729 243818 490763
rect 244026 490729 244094 490763
rect 244302 490729 244370 490763
rect 244578 490729 244646 490763
rect 244854 490729 244922 490763
rect 245130 490729 245198 490763
rect 245406 490729 245474 490763
rect 245682 490729 245750 490763
rect 245958 490729 246026 490763
rect 246234 490729 246302 490763
rect 246510 490729 246578 490763
rect 323893 372197 323961 372231
rect 324169 372197 324237 372231
rect 324445 372197 324513 372231
rect 324721 372197 324789 372231
rect 324997 372197 325065 372231
rect 325273 372197 325341 372231
rect 325549 372197 325617 372231
rect 325825 372197 325893 372231
rect 326101 372197 326169 372231
rect 326377 372197 326445 372231
rect 326653 372197 326721 372231
rect 326929 372197 326997 372231
rect 327205 372197 327273 372231
rect 327481 372197 327549 372231
rect 327757 372197 327825 372231
rect 328033 372197 328101 372231
rect 328309 372197 328377 372231
rect 328585 372197 328653 372231
rect 328861 372197 328929 372231
rect 329137 372197 329205 372231
rect 329413 372197 329481 372231
rect 329689 372197 329757 372231
rect 329965 372197 330033 372231
rect 330241 372197 330309 372231
rect 330517 372197 330585 372231
rect 330793 372197 330861 372231
rect 331069 372197 331137 372231
rect 331345 372197 331413 372231
rect 331621 372197 331689 372231
rect 331897 372197 331965 372231
rect 332173 372197 332241 372231
rect 332449 372197 332517 372231
rect 332725 372197 332793 372231
rect 333001 372197 333069 372231
rect 333277 372197 333345 372231
rect 333553 372197 333621 372231
rect 333829 372197 333897 372231
rect 334105 372197 334173 372231
rect 334381 372197 334449 372231
rect 334657 372197 334725 372231
rect 334933 372197 335001 372231
rect 335209 372197 335277 372231
rect 335485 372197 335553 372231
rect 335761 372197 335829 372231
rect 336037 372197 336105 372231
rect 336313 372197 336381 372231
rect 336589 372197 336657 372231
rect 336865 372197 336933 372231
rect 337141 372197 337209 372231
rect 337417 372197 337485 372231
rect 337693 372197 337761 372231
rect 323893 372003 323961 372037
rect 324169 372003 324237 372037
rect 324445 372003 324513 372037
rect 324721 372003 324789 372037
rect 324997 372003 325065 372037
rect 325273 372003 325341 372037
rect 325549 372003 325617 372037
rect 325825 372003 325893 372037
rect 326101 372003 326169 372037
rect 326377 372003 326445 372037
rect 326653 372003 326721 372037
rect 326929 372003 326997 372037
rect 327205 372003 327273 372037
rect 327481 372003 327549 372037
rect 327757 372003 327825 372037
rect 328033 372003 328101 372037
rect 328309 372003 328377 372037
rect 328585 372003 328653 372037
rect 328861 372003 328929 372037
rect 329137 372003 329205 372037
rect 329413 372003 329481 372037
rect 329689 372003 329757 372037
rect 329965 372003 330033 372037
rect 330241 372003 330309 372037
rect 330517 372003 330585 372037
rect 330793 372003 330861 372037
rect 331069 372003 331137 372037
rect 331345 372003 331413 372037
rect 331621 372003 331689 372037
rect 331897 372003 331965 372037
rect 332173 372003 332241 372037
rect 332449 372003 332517 372037
rect 332725 372003 332793 372037
rect 333001 372003 333069 372037
rect 333277 372003 333345 372037
rect 333553 372003 333621 372037
rect 333829 372003 333897 372037
rect 334105 372003 334173 372037
rect 334381 372003 334449 372037
rect 334657 372003 334725 372037
rect 334933 372003 335001 372037
rect 335209 372003 335277 372037
rect 335485 372003 335553 372037
rect 335761 372003 335829 372037
rect 336037 372003 336105 372037
rect 336313 372003 336381 372037
rect 336589 372003 336657 372037
rect 336865 372003 336933 372037
rect 337141 372003 337209 372037
rect 337417 372003 337485 372037
rect 337693 372003 337761 372037
rect 53353 371519 53421 371553
rect 53629 371519 53697 371553
rect 53905 371519 53973 371553
rect 54181 371519 54249 371553
rect 54457 371519 54525 371553
rect 54733 371519 54801 371553
rect 55009 371519 55077 371553
rect 55285 371519 55353 371553
rect 55561 371519 55629 371553
rect 55837 371519 55905 371553
rect 56113 371519 56181 371553
rect 56389 371519 56457 371553
rect 56665 371519 56733 371553
rect 56941 371519 57009 371553
rect 57217 371519 57285 371553
rect 57493 371519 57561 371553
rect 57769 371519 57837 371553
rect 58045 371519 58113 371553
rect 58321 371519 58389 371553
rect 58597 371519 58665 371553
rect 58873 371519 58941 371553
rect 59149 371519 59217 371553
rect 59425 371519 59493 371553
rect 59701 371519 59769 371553
rect 59977 371519 60045 371553
rect 60253 371519 60321 371553
rect 60529 371519 60597 371553
rect 60805 371519 60873 371553
rect 61081 371519 61149 371553
rect 61357 371519 61425 371553
rect 61633 371519 61701 371553
rect 61909 371519 61977 371553
rect 62185 371519 62253 371553
rect 62461 371519 62529 371553
rect 62737 371519 62805 371553
rect 63013 371519 63081 371553
rect 63289 371519 63357 371553
rect 63565 371519 63633 371553
rect 63841 371519 63909 371553
rect 64117 371519 64185 371553
rect 64393 371519 64461 371553
rect 64669 371519 64737 371553
rect 64945 371519 65013 371553
rect 65221 371519 65289 371553
rect 65497 371519 65565 371553
rect 65773 371519 65841 371553
rect 66049 371519 66117 371553
rect 66325 371519 66393 371553
rect 66601 371519 66669 371553
rect 66877 371519 66945 371553
rect 67153 371519 67221 371553
rect 53353 371325 53421 371359
rect 53629 371325 53697 371359
rect 53905 371325 53973 371359
rect 54181 371325 54249 371359
rect 54457 371325 54525 371359
rect 54733 371325 54801 371359
rect 55009 371325 55077 371359
rect 55285 371325 55353 371359
rect 55561 371325 55629 371359
rect 55837 371325 55905 371359
rect 56113 371325 56181 371359
rect 56389 371325 56457 371359
rect 56665 371325 56733 371359
rect 56941 371325 57009 371359
rect 57217 371325 57285 371359
rect 57493 371325 57561 371359
rect 57769 371325 57837 371359
rect 58045 371325 58113 371359
rect 58321 371325 58389 371359
rect 58597 371325 58665 371359
rect 58873 371325 58941 371359
rect 59149 371325 59217 371359
rect 59425 371325 59493 371359
rect 59701 371325 59769 371359
rect 59977 371325 60045 371359
rect 60253 371325 60321 371359
rect 60529 371325 60597 371359
rect 60805 371325 60873 371359
rect 61081 371325 61149 371359
rect 61357 371325 61425 371359
rect 61633 371325 61701 371359
rect 61909 371325 61977 371359
rect 62185 371325 62253 371359
rect 62461 371325 62529 371359
rect 62737 371325 62805 371359
rect 63013 371325 63081 371359
rect 63289 371325 63357 371359
rect 63565 371325 63633 371359
rect 63841 371325 63909 371359
rect 64117 371325 64185 371359
rect 64393 371325 64461 371359
rect 64669 371325 64737 371359
rect 64945 371325 65013 371359
rect 65221 371325 65289 371359
rect 65497 371325 65565 371359
rect 65773 371325 65841 371359
rect 66049 371325 66117 371359
rect 66325 371325 66393 371359
rect 66601 371325 66669 371359
rect 66877 371325 66945 371359
rect 67153 371325 67221 371359
rect 143353 371519 143421 371553
rect 143629 371519 143697 371553
rect 143905 371519 143973 371553
rect 144181 371519 144249 371553
rect 144457 371519 144525 371553
rect 144733 371519 144801 371553
rect 145009 371519 145077 371553
rect 145285 371519 145353 371553
rect 145561 371519 145629 371553
rect 145837 371519 145905 371553
rect 146113 371519 146181 371553
rect 146389 371519 146457 371553
rect 146665 371519 146733 371553
rect 146941 371519 147009 371553
rect 147217 371519 147285 371553
rect 147493 371519 147561 371553
rect 147769 371519 147837 371553
rect 148045 371519 148113 371553
rect 148321 371519 148389 371553
rect 148597 371519 148665 371553
rect 148873 371519 148941 371553
rect 149149 371519 149217 371553
rect 149425 371519 149493 371553
rect 149701 371519 149769 371553
rect 149977 371519 150045 371553
rect 150253 371519 150321 371553
rect 150529 371519 150597 371553
rect 150805 371519 150873 371553
rect 151081 371519 151149 371553
rect 151357 371519 151425 371553
rect 151633 371519 151701 371553
rect 151909 371519 151977 371553
rect 152185 371519 152253 371553
rect 152461 371519 152529 371553
rect 152737 371519 152805 371553
rect 153013 371519 153081 371553
rect 153289 371519 153357 371553
rect 153565 371519 153633 371553
rect 153841 371519 153909 371553
rect 154117 371519 154185 371553
rect 154393 371519 154461 371553
rect 154669 371519 154737 371553
rect 154945 371519 155013 371553
rect 155221 371519 155289 371553
rect 155497 371519 155565 371553
rect 155773 371519 155841 371553
rect 156049 371519 156117 371553
rect 156325 371519 156393 371553
rect 156601 371519 156669 371553
rect 156877 371519 156945 371553
rect 157153 371519 157221 371553
rect 143353 371325 143421 371359
rect 143629 371325 143697 371359
rect 143905 371325 143973 371359
rect 144181 371325 144249 371359
rect 144457 371325 144525 371359
rect 144733 371325 144801 371359
rect 145009 371325 145077 371359
rect 145285 371325 145353 371359
rect 145561 371325 145629 371359
rect 145837 371325 145905 371359
rect 146113 371325 146181 371359
rect 146389 371325 146457 371359
rect 146665 371325 146733 371359
rect 146941 371325 147009 371359
rect 147217 371325 147285 371359
rect 147493 371325 147561 371359
rect 147769 371325 147837 371359
rect 148045 371325 148113 371359
rect 148321 371325 148389 371359
rect 148597 371325 148665 371359
rect 148873 371325 148941 371359
rect 149149 371325 149217 371359
rect 149425 371325 149493 371359
rect 149701 371325 149769 371359
rect 149977 371325 150045 371359
rect 150253 371325 150321 371359
rect 150529 371325 150597 371359
rect 150805 371325 150873 371359
rect 151081 371325 151149 371359
rect 151357 371325 151425 371359
rect 151633 371325 151701 371359
rect 151909 371325 151977 371359
rect 152185 371325 152253 371359
rect 152461 371325 152529 371359
rect 152737 371325 152805 371359
rect 153013 371325 153081 371359
rect 153289 371325 153357 371359
rect 153565 371325 153633 371359
rect 153841 371325 153909 371359
rect 154117 371325 154185 371359
rect 154393 371325 154461 371359
rect 154669 371325 154737 371359
rect 154945 371325 155013 371359
rect 155221 371325 155289 371359
rect 155497 371325 155565 371359
rect 155773 371325 155841 371359
rect 156049 371325 156117 371359
rect 156325 371325 156393 371359
rect 156601 371325 156669 371359
rect 156877 371325 156945 371359
rect 157153 371325 157221 371359
rect 418903 371809 418971 371843
rect 419179 371809 419247 371843
rect 419455 371809 419523 371843
rect 419731 371809 419799 371843
rect 420007 371809 420075 371843
rect 420283 371809 420351 371843
rect 420559 371809 420627 371843
rect 420835 371809 420903 371843
rect 421111 371809 421179 371843
rect 421387 371809 421455 371843
rect 418903 371615 418971 371649
rect 419179 371615 419247 371649
rect 419455 371615 419523 371649
rect 419731 371615 419799 371649
rect 420007 371615 420075 371649
rect 420283 371615 420351 371649
rect 420559 371615 420627 371649
rect 420835 371615 420903 371649
rect 421111 371615 421179 371649
rect 421387 371615 421455 371649
rect 508902 371481 508970 371515
rect 509178 371481 509246 371515
rect 509454 371481 509522 371515
rect 509730 371481 509798 371515
rect 510006 371481 510074 371515
rect 508902 371287 508970 371321
rect 509178 371287 509246 371321
rect 509454 371287 509522 371321
rect 509730 371287 509798 371321
rect 510006 371287 510074 371321
rect 232710 370923 232778 370957
rect 232986 370923 233054 370957
rect 233262 370923 233330 370957
rect 233538 370923 233606 370957
rect 233814 370923 233882 370957
rect 234090 370923 234158 370957
rect 234366 370923 234434 370957
rect 234642 370923 234710 370957
rect 234918 370923 234986 370957
rect 235194 370923 235262 370957
rect 235470 370923 235538 370957
rect 235746 370923 235814 370957
rect 236022 370923 236090 370957
rect 236298 370923 236366 370957
rect 236574 370923 236642 370957
rect 236850 370923 236918 370957
rect 237126 370923 237194 370957
rect 237402 370923 237470 370957
rect 237678 370923 237746 370957
rect 237954 370923 238022 370957
rect 238230 370923 238298 370957
rect 238506 370923 238574 370957
rect 238782 370923 238850 370957
rect 239058 370923 239126 370957
rect 239334 370923 239402 370957
rect 239610 370923 239678 370957
rect 239886 370923 239954 370957
rect 240162 370923 240230 370957
rect 240438 370923 240506 370957
rect 240714 370923 240782 370957
rect 240990 370923 241058 370957
rect 241266 370923 241334 370957
rect 241542 370923 241610 370957
rect 241818 370923 241886 370957
rect 242094 370923 242162 370957
rect 242370 370923 242438 370957
rect 242646 370923 242714 370957
rect 242922 370923 242990 370957
rect 243198 370923 243266 370957
rect 243474 370923 243542 370957
rect 243750 370923 243818 370957
rect 244026 370923 244094 370957
rect 244302 370923 244370 370957
rect 244578 370923 244646 370957
rect 244854 370923 244922 370957
rect 245130 370923 245198 370957
rect 245406 370923 245474 370957
rect 245682 370923 245750 370957
rect 245958 370923 246026 370957
rect 246234 370923 246302 370957
rect 246510 370923 246578 370957
rect 232710 370729 232778 370763
rect 232986 370729 233054 370763
rect 233262 370729 233330 370763
rect 233538 370729 233606 370763
rect 233814 370729 233882 370763
rect 234090 370729 234158 370763
rect 234366 370729 234434 370763
rect 234642 370729 234710 370763
rect 234918 370729 234986 370763
rect 235194 370729 235262 370763
rect 235470 370729 235538 370763
rect 235746 370729 235814 370763
rect 236022 370729 236090 370763
rect 236298 370729 236366 370763
rect 236574 370729 236642 370763
rect 236850 370729 236918 370763
rect 237126 370729 237194 370763
rect 237402 370729 237470 370763
rect 237678 370729 237746 370763
rect 237954 370729 238022 370763
rect 238230 370729 238298 370763
rect 238506 370729 238574 370763
rect 238782 370729 238850 370763
rect 239058 370729 239126 370763
rect 239334 370729 239402 370763
rect 239610 370729 239678 370763
rect 239886 370729 239954 370763
rect 240162 370729 240230 370763
rect 240438 370729 240506 370763
rect 240714 370729 240782 370763
rect 240990 370729 241058 370763
rect 241266 370729 241334 370763
rect 241542 370729 241610 370763
rect 241818 370729 241886 370763
rect 242094 370729 242162 370763
rect 242370 370729 242438 370763
rect 242646 370729 242714 370763
rect 242922 370729 242990 370763
rect 243198 370729 243266 370763
rect 243474 370729 243542 370763
rect 243750 370729 243818 370763
rect 244026 370729 244094 370763
rect 244302 370729 244370 370763
rect 244578 370729 244646 370763
rect 244854 370729 244922 370763
rect 245130 370729 245198 370763
rect 245406 370729 245474 370763
rect 245682 370729 245750 370763
rect 245958 370729 246026 370763
rect 246234 370729 246302 370763
rect 246510 370729 246578 370763
rect 58902 251481 58970 251515
rect 59178 251481 59246 251515
rect 59454 251481 59522 251515
rect 59730 251481 59798 251515
rect 60006 251481 60074 251515
rect 58902 251287 58970 251321
rect 59178 251287 59246 251321
rect 59454 251287 59522 251321
rect 59730 251287 59798 251321
rect 60006 251287 60074 251321
rect 148027 251605 148095 251639
rect 148303 251605 148371 251639
rect 148579 251605 148647 251639
rect 148855 251605 148923 251639
rect 149131 251605 149199 251639
rect 149407 251605 149475 251639
rect 149683 251605 149751 251639
rect 149959 251605 150027 251639
rect 150235 251605 150303 251639
rect 150511 251605 150579 251639
rect 148027 251411 148095 251445
rect 148303 251411 148371 251445
rect 148579 251411 148647 251445
rect 148855 251411 148923 251445
rect 149131 251411 149199 251445
rect 149407 251411 149475 251445
rect 149683 251411 149751 251445
rect 149959 251411 150027 251445
rect 150235 251411 150303 251445
rect 150511 251411 150579 251445
rect 234271 251805 234339 251839
rect 234547 251805 234615 251839
rect 234823 251805 234891 251839
rect 235099 251805 235167 251839
rect 235375 251805 235443 251839
rect 235651 251805 235719 251839
rect 235927 251805 235995 251839
rect 236203 251805 236271 251839
rect 236479 251805 236547 251839
rect 236755 251805 236823 251839
rect 237031 251805 237099 251839
rect 237307 251805 237375 251839
rect 237583 251805 237651 251839
rect 237859 251805 237927 251839
rect 238135 251805 238203 251839
rect 238411 251805 238479 251839
rect 238687 251805 238755 251839
rect 238963 251805 239031 251839
rect 239239 251805 239307 251839
rect 239515 251805 239583 251839
rect 239791 251805 239859 251839
rect 240067 251805 240135 251839
rect 240343 251805 240411 251839
rect 240619 251805 240687 251839
rect 240895 251805 240963 251839
rect 241171 251805 241239 251839
rect 241447 251805 241515 251839
rect 241723 251805 241791 251839
rect 241999 251805 242067 251839
rect 242275 251805 242343 251839
rect 242551 251805 242619 251839
rect 242827 251805 242895 251839
rect 243103 251805 243171 251839
rect 243379 251805 243447 251839
rect 243655 251805 243723 251839
rect 243931 251805 243999 251839
rect 244207 251805 244275 251839
rect 244483 251805 244551 251839
rect 244759 251805 244827 251839
rect 245035 251805 245103 251839
rect 245311 251805 245379 251839
rect 245587 251805 245655 251839
rect 245863 251805 245931 251839
rect 246139 251805 246207 251839
rect 246415 251805 246483 251839
rect 246691 251805 246759 251839
rect 246967 251805 247035 251839
rect 247243 251805 247311 251839
rect 247519 251805 247587 251839
rect 247795 251805 247863 251839
rect 248071 251805 248139 251839
rect 234271 251611 234339 251645
rect 234547 251611 234615 251645
rect 234823 251611 234891 251645
rect 235099 251611 235167 251645
rect 235375 251611 235443 251645
rect 235651 251611 235719 251645
rect 235927 251611 235995 251645
rect 236203 251611 236271 251645
rect 236479 251611 236547 251645
rect 236755 251611 236823 251645
rect 237031 251611 237099 251645
rect 237307 251611 237375 251645
rect 237583 251611 237651 251645
rect 237859 251611 237927 251645
rect 238135 251611 238203 251645
rect 238411 251611 238479 251645
rect 238687 251611 238755 251645
rect 238963 251611 239031 251645
rect 239239 251611 239307 251645
rect 239515 251611 239583 251645
rect 239791 251611 239859 251645
rect 240067 251611 240135 251645
rect 240343 251611 240411 251645
rect 240619 251611 240687 251645
rect 240895 251611 240963 251645
rect 241171 251611 241239 251645
rect 241447 251611 241515 251645
rect 241723 251611 241791 251645
rect 241999 251611 242067 251645
rect 242275 251611 242343 251645
rect 242551 251611 242619 251645
rect 242827 251611 242895 251645
rect 243103 251611 243171 251645
rect 243379 251611 243447 251645
rect 243655 251611 243723 251645
rect 243931 251611 243999 251645
rect 244207 251611 244275 251645
rect 244483 251611 244551 251645
rect 244759 251611 244827 251645
rect 245035 251611 245103 251645
rect 245311 251611 245379 251645
rect 245587 251611 245655 251645
rect 245863 251611 245931 251645
rect 246139 251611 246207 251645
rect 246415 251611 246483 251645
rect 246691 251611 246759 251645
rect 246967 251611 247035 251645
rect 247243 251611 247311 251645
rect 247519 251611 247587 251645
rect 247795 251611 247863 251645
rect 248071 251611 248139 251645
rect 413353 251519 413421 251553
rect 413629 251519 413697 251553
rect 413905 251519 413973 251553
rect 414181 251519 414249 251553
rect 414457 251519 414525 251553
rect 414733 251519 414801 251553
rect 415009 251519 415077 251553
rect 415285 251519 415353 251553
rect 415561 251519 415629 251553
rect 415837 251519 415905 251553
rect 416113 251519 416181 251553
rect 416389 251519 416457 251553
rect 416665 251519 416733 251553
rect 416941 251519 417009 251553
rect 417217 251519 417285 251553
rect 417493 251519 417561 251553
rect 417769 251519 417837 251553
rect 418045 251519 418113 251553
rect 418321 251519 418389 251553
rect 418597 251519 418665 251553
rect 418873 251519 418941 251553
rect 419149 251519 419217 251553
rect 419425 251519 419493 251553
rect 419701 251519 419769 251553
rect 419977 251519 420045 251553
rect 420253 251519 420321 251553
rect 420529 251519 420597 251553
rect 420805 251519 420873 251553
rect 421081 251519 421149 251553
rect 421357 251519 421425 251553
rect 421633 251519 421701 251553
rect 421909 251519 421977 251553
rect 422185 251519 422253 251553
rect 422461 251519 422529 251553
rect 422737 251519 422805 251553
rect 423013 251519 423081 251553
rect 423289 251519 423357 251553
rect 423565 251519 423633 251553
rect 423841 251519 423909 251553
rect 424117 251519 424185 251553
rect 424393 251519 424461 251553
rect 424669 251519 424737 251553
rect 424945 251519 425013 251553
rect 425221 251519 425289 251553
rect 425497 251519 425565 251553
rect 425773 251519 425841 251553
rect 426049 251519 426117 251553
rect 426325 251519 426393 251553
rect 426601 251519 426669 251553
rect 426877 251519 426945 251553
rect 427153 251519 427221 251553
rect 413353 251325 413421 251359
rect 413629 251325 413697 251359
rect 413905 251325 413973 251359
rect 414181 251325 414249 251359
rect 414457 251325 414525 251359
rect 414733 251325 414801 251359
rect 415009 251325 415077 251359
rect 415285 251325 415353 251359
rect 415561 251325 415629 251359
rect 415837 251325 415905 251359
rect 416113 251325 416181 251359
rect 416389 251325 416457 251359
rect 416665 251325 416733 251359
rect 416941 251325 417009 251359
rect 417217 251325 417285 251359
rect 417493 251325 417561 251359
rect 417769 251325 417837 251359
rect 418045 251325 418113 251359
rect 418321 251325 418389 251359
rect 418597 251325 418665 251359
rect 418873 251325 418941 251359
rect 419149 251325 419217 251359
rect 419425 251325 419493 251359
rect 419701 251325 419769 251359
rect 419977 251325 420045 251359
rect 420253 251325 420321 251359
rect 420529 251325 420597 251359
rect 420805 251325 420873 251359
rect 421081 251325 421149 251359
rect 421357 251325 421425 251359
rect 421633 251325 421701 251359
rect 421909 251325 421977 251359
rect 422185 251325 422253 251359
rect 422461 251325 422529 251359
rect 422737 251325 422805 251359
rect 423013 251325 423081 251359
rect 423289 251325 423357 251359
rect 423565 251325 423633 251359
rect 423841 251325 423909 251359
rect 424117 251325 424185 251359
rect 424393 251325 424461 251359
rect 424669 251325 424737 251359
rect 424945 251325 425013 251359
rect 425221 251325 425289 251359
rect 425497 251325 425565 251359
rect 425773 251325 425841 251359
rect 426049 251325 426117 251359
rect 426325 251325 426393 251359
rect 426601 251325 426669 251359
rect 426877 251325 426945 251359
rect 427153 251325 427221 251359
rect 503353 251519 503421 251553
rect 503629 251519 503697 251553
rect 503905 251519 503973 251553
rect 504181 251519 504249 251553
rect 504457 251519 504525 251553
rect 504733 251519 504801 251553
rect 505009 251519 505077 251553
rect 505285 251519 505353 251553
rect 505561 251519 505629 251553
rect 505837 251519 505905 251553
rect 506113 251519 506181 251553
rect 506389 251519 506457 251553
rect 506665 251519 506733 251553
rect 506941 251519 507009 251553
rect 507217 251519 507285 251553
rect 507493 251519 507561 251553
rect 507769 251519 507837 251553
rect 508045 251519 508113 251553
rect 508321 251519 508389 251553
rect 508597 251519 508665 251553
rect 508873 251519 508941 251553
rect 509149 251519 509217 251553
rect 509425 251519 509493 251553
rect 509701 251519 509769 251553
rect 509977 251519 510045 251553
rect 510253 251519 510321 251553
rect 510529 251519 510597 251553
rect 510805 251519 510873 251553
rect 511081 251519 511149 251553
rect 511357 251519 511425 251553
rect 511633 251519 511701 251553
rect 511909 251519 511977 251553
rect 512185 251519 512253 251553
rect 512461 251519 512529 251553
rect 512737 251519 512805 251553
rect 513013 251519 513081 251553
rect 513289 251519 513357 251553
rect 513565 251519 513633 251553
rect 513841 251519 513909 251553
rect 514117 251519 514185 251553
rect 514393 251519 514461 251553
rect 514669 251519 514737 251553
rect 514945 251519 515013 251553
rect 515221 251519 515289 251553
rect 515497 251519 515565 251553
rect 515773 251519 515841 251553
rect 516049 251519 516117 251553
rect 516325 251519 516393 251553
rect 516601 251519 516669 251553
rect 516877 251519 516945 251553
rect 517153 251519 517221 251553
rect 503353 251325 503421 251359
rect 503629 251325 503697 251359
rect 503905 251325 503973 251359
rect 504181 251325 504249 251359
rect 504457 251325 504525 251359
rect 504733 251325 504801 251359
rect 505009 251325 505077 251359
rect 505285 251325 505353 251359
rect 505561 251325 505629 251359
rect 505837 251325 505905 251359
rect 506113 251325 506181 251359
rect 506389 251325 506457 251359
rect 506665 251325 506733 251359
rect 506941 251325 507009 251359
rect 507217 251325 507285 251359
rect 507493 251325 507561 251359
rect 507769 251325 507837 251359
rect 508045 251325 508113 251359
rect 508321 251325 508389 251359
rect 508597 251325 508665 251359
rect 508873 251325 508941 251359
rect 509149 251325 509217 251359
rect 509425 251325 509493 251359
rect 509701 251325 509769 251359
rect 509977 251325 510045 251359
rect 510253 251325 510321 251359
rect 510529 251325 510597 251359
rect 510805 251325 510873 251359
rect 511081 251325 511149 251359
rect 511357 251325 511425 251359
rect 511633 251325 511701 251359
rect 511909 251325 511977 251359
rect 512185 251325 512253 251359
rect 512461 251325 512529 251359
rect 512737 251325 512805 251359
rect 513013 251325 513081 251359
rect 513289 251325 513357 251359
rect 513565 251325 513633 251359
rect 513841 251325 513909 251359
rect 514117 251325 514185 251359
rect 514393 251325 514461 251359
rect 514669 251325 514737 251359
rect 514945 251325 515013 251359
rect 515221 251325 515289 251359
rect 515497 251325 515565 251359
rect 515773 251325 515841 251359
rect 516049 251325 516117 251359
rect 516325 251325 516393 251359
rect 516601 251325 516669 251359
rect 516877 251325 516945 251359
rect 517153 251325 517221 251359
rect 322710 250923 322778 250957
rect 322986 250923 323054 250957
rect 323262 250923 323330 250957
rect 323538 250923 323606 250957
rect 323814 250923 323882 250957
rect 324090 250923 324158 250957
rect 324366 250923 324434 250957
rect 324642 250923 324710 250957
rect 324918 250923 324986 250957
rect 325194 250923 325262 250957
rect 325470 250923 325538 250957
rect 325746 250923 325814 250957
rect 326022 250923 326090 250957
rect 326298 250923 326366 250957
rect 326574 250923 326642 250957
rect 326850 250923 326918 250957
rect 327126 250923 327194 250957
rect 327402 250923 327470 250957
rect 327678 250923 327746 250957
rect 327954 250923 328022 250957
rect 328230 250923 328298 250957
rect 328506 250923 328574 250957
rect 328782 250923 328850 250957
rect 329058 250923 329126 250957
rect 329334 250923 329402 250957
rect 329610 250923 329678 250957
rect 329886 250923 329954 250957
rect 330162 250923 330230 250957
rect 330438 250923 330506 250957
rect 330714 250923 330782 250957
rect 330990 250923 331058 250957
rect 331266 250923 331334 250957
rect 331542 250923 331610 250957
rect 331818 250923 331886 250957
rect 332094 250923 332162 250957
rect 332370 250923 332438 250957
rect 332646 250923 332714 250957
rect 332922 250923 332990 250957
rect 333198 250923 333266 250957
rect 333474 250923 333542 250957
rect 333750 250923 333818 250957
rect 334026 250923 334094 250957
rect 334302 250923 334370 250957
rect 334578 250923 334646 250957
rect 334854 250923 334922 250957
rect 335130 250923 335198 250957
rect 335406 250923 335474 250957
rect 335682 250923 335750 250957
rect 335958 250923 336026 250957
rect 336234 250923 336302 250957
rect 336510 250923 336578 250957
rect 322710 250729 322778 250763
rect 322986 250729 323054 250763
rect 323262 250729 323330 250763
rect 323538 250729 323606 250763
rect 323814 250729 323882 250763
rect 324090 250729 324158 250763
rect 324366 250729 324434 250763
rect 324642 250729 324710 250763
rect 324918 250729 324986 250763
rect 325194 250729 325262 250763
rect 325470 250729 325538 250763
rect 325746 250729 325814 250763
rect 326022 250729 326090 250763
rect 326298 250729 326366 250763
rect 326574 250729 326642 250763
rect 326850 250729 326918 250763
rect 327126 250729 327194 250763
rect 327402 250729 327470 250763
rect 327678 250729 327746 250763
rect 327954 250729 328022 250763
rect 328230 250729 328298 250763
rect 328506 250729 328574 250763
rect 328782 250729 328850 250763
rect 329058 250729 329126 250763
rect 329334 250729 329402 250763
rect 329610 250729 329678 250763
rect 329886 250729 329954 250763
rect 330162 250729 330230 250763
rect 330438 250729 330506 250763
rect 330714 250729 330782 250763
rect 330990 250729 331058 250763
rect 331266 250729 331334 250763
rect 331542 250729 331610 250763
rect 331818 250729 331886 250763
rect 332094 250729 332162 250763
rect 332370 250729 332438 250763
rect 332646 250729 332714 250763
rect 332922 250729 332990 250763
rect 333198 250729 333266 250763
rect 333474 250729 333542 250763
rect 333750 250729 333818 250763
rect 334026 250729 334094 250763
rect 334302 250729 334370 250763
rect 334578 250729 334646 250763
rect 334854 250729 334922 250763
rect 335130 250729 335198 250763
rect 335406 250729 335474 250763
rect 335682 250729 335750 250763
rect 335958 250729 336026 250763
rect 336234 250729 336302 250763
rect 336510 250729 336578 250763
rect 59339 145993 59373 146027
rect 59339 145665 59373 145699
rect 149537 145589 149605 145623
rect 149537 145261 149605 145295
rect 239356 146022 239390 146056
rect 239356 145712 239390 145746
rect 329339 145993 329373 146027
rect 329339 145665 329373 145699
rect 419537 145589 419605 145623
rect 419537 145261 419605 145295
rect 509356 146022 509390 146056
rect 509356 145712 509390 145746
rect 59356 56022 59390 56056
rect 59356 55712 59390 55746
rect 149627 56021 149695 56055
rect 149627 55711 149695 55745
rect 239637 55731 239705 55765
rect 239637 55421 239705 55455
rect 329356 56022 329390 56056
rect 329356 55712 329390 55746
rect 419627 56021 419695 56055
rect 419627 55711 419695 55745
rect 509637 55731 509705 55765
rect 509637 55421 509705 55455
<< locali >>
rect 329316 657986 329350 658002
rect 329142 657946 329158 657980
rect 329192 657946 329208 657980
rect 329114 657896 329148 657912
rect 329114 657704 329148 657720
rect 329202 657896 329236 657912
rect 329202 657704 329236 657720
rect 329142 657636 329158 657670
rect 329192 657636 329208 657670
rect 509316 657986 509350 658002
rect 509142 657946 509158 657980
rect 509192 657946 509208 657980
rect 509114 657896 509148 657912
rect 509114 657704 509148 657720
rect 509202 657896 509236 657912
rect 509202 657704 509236 657720
rect 509142 657636 509158 657670
rect 509192 657636 509208 657670
rect 329316 657614 329350 657630
rect 509316 657614 509350 657630
rect 419569 657589 419603 657605
rect 419323 657513 419339 657547
rect 419407 657513 419423 657547
rect 419277 657454 419311 657470
rect 419277 657262 419311 657278
rect 419435 657454 419469 657470
rect 419435 657262 419469 657278
rect 419323 657185 419339 657219
rect 419407 657185 419423 657219
rect 419569 657127 419603 657143
rect 59857 656097 59891 656113
rect 59611 656021 59627 656055
rect 59695 656021 59711 656055
rect 59565 655971 59599 655987
rect 59565 655779 59599 655795
rect 59723 655971 59757 655987
rect 59723 655779 59757 655795
rect 59611 655711 59627 655745
rect 59695 655711 59711 655745
rect 149514 656062 149548 656078
rect 149340 656022 149356 656056
rect 149390 656022 149406 656056
rect 149312 655972 149346 655988
rect 149312 655780 149346 655796
rect 149400 655972 149434 655988
rect 149400 655780 149434 655796
rect 149340 655712 149356 655746
rect 149390 655712 149406 655746
rect 239497 656033 239531 656049
rect 239323 655993 239339 656027
rect 239373 655993 239389 656027
rect 239295 655934 239329 655950
rect 239295 655742 239329 655758
rect 239383 655934 239417 655950
rect 239383 655742 239417 655758
rect 149514 655690 149548 655706
rect 59857 655653 59891 655669
rect 239323 655665 239339 655699
rect 239373 655665 239389 655699
rect 239497 655643 239531 655659
rect 419659 583021 419693 583037
rect 419413 582945 419429 582979
rect 419497 582945 419513 582979
rect 419367 582895 419401 582911
rect 419367 582703 419401 582719
rect 419525 582895 419559 582911
rect 419525 582703 419559 582719
rect 419413 582635 419429 582669
rect 419497 582635 419513 582669
rect 509669 582731 509703 582747
rect 509423 582655 509439 582689
rect 509507 582655 509523 582689
rect 419659 582577 419693 582593
rect 509377 582605 509411 582621
rect 509377 582413 509411 582429
rect 509535 582605 509569 582621
rect 509535 582413 509569 582429
rect 509423 582345 509439 582379
rect 509507 582345 509523 582379
rect 509669 582287 509703 582303
rect 59857 581097 59891 581113
rect 59611 581021 59627 581055
rect 59695 581021 59711 581055
rect 59565 580971 59599 580987
rect 59565 580779 59599 580795
rect 59723 580971 59757 580987
rect 59723 580779 59757 580795
rect 59611 580711 59627 580745
rect 59695 580711 59711 580745
rect 239514 581062 239548 581078
rect 239340 581022 239356 581056
rect 239390 581022 239406 581056
rect 239312 580972 239346 580988
rect 149867 580807 149901 580823
rect 149621 580731 149637 580765
rect 149705 580731 149721 580765
rect 59857 580653 59891 580669
rect 149575 580681 149609 580697
rect 149575 580489 149609 580505
rect 149733 580681 149767 580697
rect 149733 580489 149767 580505
rect 149621 580421 149637 580455
rect 149705 580421 149721 580455
rect 239312 580780 239346 580796
rect 239400 580972 239434 580988
rect 239400 580780 239434 580796
rect 239340 580712 239356 580746
rect 239390 580712 239406 580746
rect 239514 580690 239548 580706
rect 329767 580665 329801 580681
rect 329521 580589 329537 580623
rect 329605 580589 329621 580623
rect 149867 580363 149901 580379
rect 329475 580530 329509 580546
rect 329475 580338 329509 580354
rect 329633 580530 329667 580546
rect 329633 580338 329667 580354
rect 329521 580261 329537 580295
rect 329605 580261 329621 580295
rect 329767 580203 329801 580219
rect 323888 492598 323968 492608
rect 323888 492556 323904 492598
rect 323958 492556 323968 492598
rect 323888 492231 323968 492556
rect 324161 492488 338373 492515
rect 324160 492417 338373 492488
rect 324160 492231 324258 492417
rect 324436 492231 324534 492417
rect 324710 492231 324808 492417
rect 324988 492231 325086 492417
rect 325260 492231 325358 492417
rect 325538 492231 325636 492417
rect 325816 492231 325914 492417
rect 326094 492231 326192 492417
rect 326368 492231 326466 492417
rect 326644 492231 326742 492417
rect 326920 492231 327018 492417
rect 327198 492231 327296 492417
rect 327474 492231 327572 492417
rect 327746 492231 327844 492417
rect 328024 492231 328122 492417
rect 328296 492231 328394 492417
rect 328574 492231 328672 492417
rect 328850 492231 328948 492417
rect 323877 492197 323893 492231
rect 323961 492197 323977 492231
rect 324153 492197 324169 492231
rect 324237 492206 324258 492231
rect 324237 492197 324253 492206
rect 324429 492197 324445 492231
rect 324513 492208 324534 492231
rect 324513 492197 324529 492208
rect 324705 492197 324721 492231
rect 324789 492204 324808 492231
rect 324789 492197 324805 492204
rect 324981 492197 324997 492231
rect 325065 492204 325086 492231
rect 325065 492197 325081 492204
rect 325257 492197 325273 492231
rect 325341 492206 325358 492231
rect 325341 492197 325357 492206
rect 325533 492197 325549 492231
rect 325617 492204 325636 492231
rect 325617 492197 325633 492204
rect 325809 492197 325825 492231
rect 325893 492204 325914 492231
rect 325893 492197 325909 492204
rect 326085 492197 326101 492231
rect 326169 492208 326192 492231
rect 326169 492197 326185 492208
rect 326361 492197 326377 492231
rect 326445 492204 326466 492231
rect 326445 492197 326461 492204
rect 326637 492197 326653 492231
rect 326721 492208 326742 492231
rect 326721 492197 326737 492208
rect 326913 492197 326929 492231
rect 326997 492208 327018 492231
rect 326997 492197 327013 492208
rect 327189 492197 327205 492231
rect 327273 492210 327296 492231
rect 327273 492197 327289 492210
rect 327465 492197 327481 492231
rect 327549 492200 327572 492231
rect 327549 492197 327565 492200
rect 327741 492197 327757 492231
rect 327825 492204 327844 492231
rect 327825 492197 327841 492204
rect 328017 492197 328033 492231
rect 328101 492204 328122 492231
rect 328101 492197 328117 492204
rect 328293 492197 328309 492231
rect 328377 492197 328394 492231
rect 328569 492197 328585 492231
rect 328653 492204 328672 492231
rect 328653 492197 328669 492204
rect 328845 492197 328861 492231
rect 328929 492204 328948 492231
rect 329120 492231 329218 492417
rect 329406 492231 329504 492417
rect 329678 492231 329776 492417
rect 329958 492231 330056 492417
rect 330232 492231 330330 492417
rect 330508 492231 330606 492417
rect 330784 492231 330882 492417
rect 331060 492231 331158 492417
rect 331336 492231 331434 492417
rect 331612 492231 331710 492417
rect 331888 492231 331986 492417
rect 332164 492231 332262 492417
rect 332442 492231 332540 492417
rect 332718 492231 332816 492417
rect 332990 492231 333088 492417
rect 333268 492231 333366 492417
rect 333544 492231 333642 492417
rect 333822 492231 333920 492417
rect 334096 492231 334194 492417
rect 334372 492231 334470 492417
rect 334650 492231 334748 492417
rect 334926 492231 335024 492417
rect 335202 492231 335300 492417
rect 335478 492231 335576 492417
rect 335754 492231 335852 492417
rect 336028 492231 336126 492417
rect 336308 492231 336406 492417
rect 336584 492231 336682 492417
rect 336856 492231 336954 492417
rect 337132 492231 337230 492417
rect 337402 492231 337500 492417
rect 337694 492231 337792 492417
rect 328929 492197 328945 492204
rect 329120 492202 329137 492231
rect 329121 492197 329137 492202
rect 329205 492197 329221 492231
rect 329397 492197 329413 492231
rect 329481 492200 329504 492231
rect 329481 492197 329497 492200
rect 329673 492197 329689 492231
rect 329757 492200 329776 492231
rect 329757 492197 329773 492200
rect 329949 492197 329965 492231
rect 330033 492200 330056 492231
rect 330033 492197 330049 492200
rect 330225 492197 330241 492231
rect 330309 492200 330330 492231
rect 330309 492197 330325 492200
rect 330501 492197 330517 492231
rect 330585 492202 330606 492231
rect 330585 492197 330601 492202
rect 330777 492197 330793 492231
rect 330861 492200 330882 492231
rect 330861 492197 330877 492200
rect 331053 492197 331069 492231
rect 331137 492202 331158 492231
rect 331137 492197 331153 492202
rect 331329 492197 331345 492231
rect 331413 492202 331434 492231
rect 331413 492197 331429 492202
rect 331605 492197 331621 492231
rect 331689 492204 331710 492231
rect 331689 492197 331705 492204
rect 331881 492197 331897 492231
rect 331965 492202 331986 492231
rect 331965 492197 331981 492202
rect 332157 492197 332173 492231
rect 332241 492202 332262 492231
rect 332241 492197 332257 492202
rect 332433 492197 332449 492231
rect 332517 492202 332540 492231
rect 332517 492197 332533 492202
rect 332709 492197 332725 492231
rect 332793 492202 332816 492231
rect 332793 492197 332809 492202
rect 332985 492197 333001 492231
rect 333069 492200 333088 492231
rect 333069 492197 333085 492200
rect 333261 492197 333277 492231
rect 333345 492200 333366 492231
rect 333345 492197 333361 492200
rect 333537 492197 333553 492231
rect 333621 492204 333642 492231
rect 333621 492197 333637 492204
rect 333813 492197 333829 492231
rect 333897 492206 333920 492231
rect 333897 492197 333913 492206
rect 334089 492197 334105 492231
rect 334173 492202 334194 492231
rect 334173 492197 334189 492202
rect 334365 492197 334381 492231
rect 334449 492206 334470 492231
rect 334449 492197 334465 492206
rect 334641 492197 334657 492231
rect 334725 492206 334748 492231
rect 334725 492197 334741 492206
rect 334917 492197 334933 492231
rect 335001 492208 335024 492231
rect 335001 492197 335017 492208
rect 335193 492197 335209 492231
rect 335277 492204 335300 492231
rect 335277 492197 335293 492204
rect 335469 492197 335485 492231
rect 335553 492206 335576 492231
rect 335553 492197 335569 492206
rect 335745 492197 335761 492231
rect 335829 492206 335852 492231
rect 335829 492197 335845 492206
rect 336021 492197 336037 492231
rect 336105 492208 336126 492231
rect 336105 492197 336121 492208
rect 336297 492197 336313 492231
rect 336381 492208 336406 492231
rect 336381 492197 336397 492208
rect 336573 492197 336589 492231
rect 336657 492208 336682 492231
rect 336657 492197 336673 492208
rect 336849 492197 336865 492231
rect 336933 492208 336954 492231
rect 336933 492197 336949 492208
rect 337125 492197 337141 492231
rect 337209 492198 337230 492231
rect 337209 492197 337225 492198
rect 337401 492197 337417 492231
rect 337485 492197 337501 492231
rect 337677 492197 337693 492231
rect 337761 492198 337792 492231
rect 337923 492273 337957 492289
rect 337761 492197 337777 492198
rect 323888 492192 323968 492197
rect 328296 492196 328394 492197
rect 337402 492196 337500 492197
rect 323831 492147 323865 492163
rect 323831 492071 323865 492087
rect 323989 492147 324023 492163
rect 323989 492071 324023 492087
rect 324107 492147 324141 492163
rect 324107 492071 324141 492087
rect 324265 492147 324299 492163
rect 324265 492071 324299 492087
rect 324383 492147 324417 492163
rect 324383 492071 324417 492087
rect 324541 492147 324575 492163
rect 324541 492071 324575 492087
rect 324659 492147 324693 492163
rect 324659 492071 324693 492087
rect 324817 492147 324851 492163
rect 324817 492071 324851 492087
rect 324935 492147 324969 492163
rect 324935 492071 324969 492087
rect 325093 492147 325127 492163
rect 325093 492071 325127 492087
rect 325211 492147 325245 492163
rect 325211 492071 325245 492087
rect 325369 492147 325403 492163
rect 325369 492071 325403 492087
rect 325487 492147 325521 492163
rect 325487 492071 325521 492087
rect 325645 492147 325679 492163
rect 325645 492071 325679 492087
rect 325763 492147 325797 492163
rect 325763 492071 325797 492087
rect 325921 492147 325955 492163
rect 325921 492071 325955 492087
rect 326039 492147 326073 492163
rect 326039 492071 326073 492087
rect 326197 492147 326231 492163
rect 326197 492071 326231 492087
rect 326315 492147 326349 492163
rect 326315 492071 326349 492087
rect 326473 492147 326507 492163
rect 326473 492071 326507 492087
rect 326591 492147 326625 492163
rect 326591 492071 326625 492087
rect 326749 492147 326783 492163
rect 326749 492071 326783 492087
rect 326867 492147 326901 492163
rect 326867 492071 326901 492087
rect 327025 492147 327059 492163
rect 327025 492071 327059 492087
rect 327143 492147 327177 492163
rect 327143 492071 327177 492087
rect 327301 492147 327335 492163
rect 327301 492071 327335 492087
rect 327419 492147 327453 492163
rect 327419 492071 327453 492087
rect 327577 492147 327611 492163
rect 327577 492071 327611 492087
rect 327695 492147 327729 492163
rect 327695 492071 327729 492087
rect 327853 492147 327887 492163
rect 327853 492071 327887 492087
rect 327971 492147 328005 492163
rect 327971 492071 328005 492087
rect 328129 492147 328163 492163
rect 328129 492071 328163 492087
rect 328247 492147 328281 492163
rect 328247 492071 328281 492087
rect 328405 492147 328439 492163
rect 328405 492071 328439 492087
rect 328523 492147 328557 492163
rect 328523 492071 328557 492087
rect 328681 492147 328715 492163
rect 328681 492071 328715 492087
rect 328799 492147 328833 492163
rect 328799 492071 328833 492087
rect 328957 492147 328991 492163
rect 328957 492071 328991 492087
rect 329075 492147 329109 492163
rect 329075 492071 329109 492087
rect 329233 492147 329267 492163
rect 329233 492071 329267 492087
rect 329351 492147 329385 492163
rect 329351 492071 329385 492087
rect 329509 492147 329543 492163
rect 329509 492071 329543 492087
rect 329627 492147 329661 492163
rect 329627 492071 329661 492087
rect 329785 492147 329819 492163
rect 329785 492071 329819 492087
rect 329903 492147 329937 492163
rect 329903 492071 329937 492087
rect 330061 492147 330095 492163
rect 330061 492071 330095 492087
rect 330179 492147 330213 492163
rect 330179 492071 330213 492087
rect 330337 492147 330371 492163
rect 330337 492071 330371 492087
rect 330455 492147 330489 492163
rect 330455 492071 330489 492087
rect 330613 492147 330647 492163
rect 330613 492071 330647 492087
rect 330731 492147 330765 492163
rect 330731 492071 330765 492087
rect 330889 492147 330923 492163
rect 330889 492071 330923 492087
rect 331007 492147 331041 492163
rect 331007 492071 331041 492087
rect 331165 492147 331199 492163
rect 331165 492071 331199 492087
rect 331283 492147 331317 492163
rect 331283 492071 331317 492087
rect 331441 492147 331475 492163
rect 331441 492071 331475 492087
rect 331559 492147 331593 492163
rect 331559 492071 331593 492087
rect 331717 492147 331751 492163
rect 331717 492071 331751 492087
rect 331835 492147 331869 492163
rect 331835 492071 331869 492087
rect 331993 492147 332027 492163
rect 331993 492071 332027 492087
rect 332111 492147 332145 492163
rect 332111 492071 332145 492087
rect 332269 492147 332303 492163
rect 332269 492071 332303 492087
rect 332387 492147 332421 492163
rect 332387 492071 332421 492087
rect 332545 492147 332579 492163
rect 332545 492071 332579 492087
rect 332663 492147 332697 492163
rect 332663 492071 332697 492087
rect 332821 492147 332855 492163
rect 332821 492071 332855 492087
rect 332939 492147 332973 492163
rect 332939 492071 332973 492087
rect 333097 492147 333131 492163
rect 333097 492071 333131 492087
rect 333215 492147 333249 492163
rect 333215 492071 333249 492087
rect 333373 492147 333407 492163
rect 333373 492071 333407 492087
rect 333491 492147 333525 492163
rect 333491 492071 333525 492087
rect 333649 492147 333683 492163
rect 333649 492071 333683 492087
rect 333767 492147 333801 492163
rect 333767 492071 333801 492087
rect 333925 492147 333959 492163
rect 333925 492071 333959 492087
rect 334043 492147 334077 492163
rect 334043 492071 334077 492087
rect 334201 492147 334235 492163
rect 334201 492071 334235 492087
rect 334319 492147 334353 492163
rect 334319 492071 334353 492087
rect 334477 492147 334511 492163
rect 334477 492071 334511 492087
rect 334595 492147 334629 492163
rect 334595 492071 334629 492087
rect 334753 492147 334787 492163
rect 334753 492071 334787 492087
rect 334871 492147 334905 492163
rect 334871 492071 334905 492087
rect 335029 492147 335063 492163
rect 335029 492071 335063 492087
rect 335147 492147 335181 492163
rect 335147 492071 335181 492087
rect 335305 492147 335339 492163
rect 335305 492071 335339 492087
rect 335423 492147 335457 492163
rect 335423 492071 335457 492087
rect 335581 492147 335615 492163
rect 335581 492071 335615 492087
rect 335699 492147 335733 492163
rect 335699 492071 335733 492087
rect 335857 492147 335891 492163
rect 335857 492071 335891 492087
rect 335975 492147 336009 492163
rect 335975 492071 336009 492087
rect 336133 492147 336167 492163
rect 336133 492071 336167 492087
rect 336251 492147 336285 492163
rect 336251 492071 336285 492087
rect 336409 492147 336443 492163
rect 336409 492071 336443 492087
rect 336527 492147 336561 492163
rect 336527 492071 336561 492087
rect 336685 492147 336719 492163
rect 336685 492071 336719 492087
rect 336803 492147 336837 492163
rect 336803 492071 336837 492087
rect 336961 492147 336995 492163
rect 336961 492071 336995 492087
rect 337079 492147 337113 492163
rect 337079 492071 337113 492087
rect 337237 492147 337271 492163
rect 337237 492071 337271 492087
rect 337355 492147 337389 492163
rect 337355 492071 337389 492087
rect 337513 492147 337547 492163
rect 337513 492071 337547 492087
rect 337631 492147 337665 492163
rect 337631 492071 337665 492087
rect 337789 492147 337823 492163
rect 337789 492071 337823 492087
rect 323888 492037 323968 492040
rect 323877 492003 323893 492037
rect 323961 492003 323977 492037
rect 324153 492003 324169 492037
rect 324237 492003 324253 492037
rect 324429 492032 324445 492037
rect 324426 492003 324445 492032
rect 324513 492003 324529 492037
rect 324705 492028 324721 492037
rect 324702 492003 324721 492028
rect 324789 492003 324805 492037
rect 324981 492022 324997 492037
rect 324980 492003 324997 492022
rect 325065 492003 325081 492037
rect 325257 492018 325273 492037
rect 325256 492003 325273 492018
rect 325341 492003 325357 492037
rect 325533 492020 325549 492037
rect 325530 492003 325549 492020
rect 325617 492003 325633 492037
rect 325809 492018 325825 492037
rect 325808 492003 325825 492018
rect 325893 492003 325909 492037
rect 326085 492003 326101 492037
rect 326169 492003 326185 492037
rect 326361 492018 326377 492037
rect 326360 492003 326377 492018
rect 326445 492003 326461 492037
rect 326637 492003 326653 492037
rect 326721 492003 326737 492037
rect 326913 492028 326929 492037
rect 326910 492003 326929 492028
rect 326997 492003 327013 492037
rect 327189 492028 327205 492037
rect 327186 492003 327205 492028
rect 327273 492003 327289 492037
rect 327465 492003 327481 492037
rect 327549 492003 327565 492037
rect 327741 492022 327757 492037
rect 327734 492003 327757 492022
rect 327825 492003 327841 492037
rect 328017 492003 328033 492037
rect 328101 492003 328117 492037
rect 328293 492022 328309 492037
rect 328292 492003 328309 492022
rect 328377 492003 328393 492037
rect 328569 492018 328585 492037
rect 328568 492003 328585 492018
rect 328653 492003 328669 492037
rect 328845 492026 328861 492037
rect 328842 492003 328861 492026
rect 328929 492003 328945 492037
rect 329121 492018 329137 492037
rect 329120 492003 329137 492018
rect 329205 492003 329221 492037
rect 329397 492020 329413 492037
rect 329390 492003 329413 492020
rect 329481 492003 329497 492037
rect 329673 492026 329689 492037
rect 329666 492003 329689 492026
rect 329757 492003 329773 492037
rect 329949 492032 329965 492037
rect 329948 492003 329965 492032
rect 330033 492003 330049 492037
rect 330225 492028 330241 492037
rect 330224 492003 330241 492028
rect 330309 492003 330325 492037
rect 330501 492028 330517 492037
rect 330498 492003 330517 492028
rect 330585 492003 330601 492037
rect 330777 492028 330793 492037
rect 330770 492003 330793 492028
rect 330861 492003 330877 492037
rect 331053 492028 331069 492037
rect 331052 492003 331069 492028
rect 331137 492003 331153 492037
rect 331329 492003 331345 492037
rect 331413 492003 331429 492037
rect 331605 492022 331621 492037
rect 331604 492003 331621 492022
rect 331689 492003 331705 492037
rect 331881 492003 331897 492037
rect 331965 492003 331981 492037
rect 332157 492003 332173 492037
rect 332241 492003 332257 492037
rect 332433 492014 332449 492037
rect 332426 492003 332449 492014
rect 332517 492003 332533 492037
rect 332709 492010 332725 492037
rect 332708 492003 332725 492010
rect 332793 492003 332809 492037
rect 332985 492003 333001 492037
rect 333069 492003 333085 492037
rect 333261 492010 333277 492037
rect 333260 492003 333277 492010
rect 333345 492003 333361 492037
rect 333537 492010 333553 492037
rect 333536 492003 333553 492010
rect 333621 492003 333637 492037
rect 333813 492026 333829 492037
rect 333806 492003 333829 492026
rect 333897 492003 333913 492037
rect 334089 492018 334105 492037
rect 334084 492003 334105 492018
rect 334173 492003 334189 492037
rect 334365 492003 334381 492037
rect 334449 492003 334465 492037
rect 334641 492003 334657 492037
rect 334725 492018 334741 492037
rect 334917 492022 334933 492037
rect 334725 492003 334746 492018
rect 58580 491988 61459 491999
rect 58580 491957 61460 491988
rect 58580 491514 58622 491957
rect 58900 491952 61460 491957
rect 58900 491843 58978 491952
rect 59176 491843 59254 491952
rect 59454 491843 59532 491952
rect 59726 491843 59804 491952
rect 60008 491843 60086 491850
rect 60280 491843 60358 491952
rect 60556 491843 60634 491952
rect 60830 491843 60908 491952
rect 61108 491843 61186 491952
rect 61382 491843 61460 491952
rect 61617 491885 61651 491901
rect 58887 491809 58903 491843
rect 58971 491809 58987 491843
rect 59163 491809 59179 491843
rect 59247 491809 59263 491843
rect 59439 491809 59455 491843
rect 59523 491809 59539 491843
rect 59715 491809 59731 491843
rect 59799 491809 59815 491843
rect 59991 491809 60007 491843
rect 60075 491809 60091 491843
rect 60267 491809 60283 491843
rect 60351 491809 60367 491843
rect 60543 491809 60559 491843
rect 60627 491809 60643 491843
rect 60819 491809 60835 491843
rect 60903 491809 60919 491843
rect 61095 491809 61111 491843
rect 61179 491809 61195 491843
rect 61371 491809 61387 491843
rect 61455 491809 61471 491843
rect 58900 491808 58978 491809
rect 59176 491806 59254 491809
rect 59454 491808 59532 491809
rect 59726 491808 59804 491809
rect 60008 491808 60086 491809
rect 60280 491808 60358 491809
rect 60556 491806 60634 491809
rect 60830 491806 60908 491809
rect 61108 491808 61186 491809
rect 61382 491806 61460 491809
rect 58841 491759 58875 491775
rect 58841 491683 58875 491699
rect 58999 491759 59033 491775
rect 58999 491683 59033 491699
rect 59117 491759 59151 491775
rect 59117 491683 59151 491699
rect 59275 491759 59309 491775
rect 59275 491683 59309 491699
rect 59393 491759 59427 491775
rect 59393 491683 59427 491699
rect 59551 491759 59585 491775
rect 59551 491683 59585 491699
rect 59669 491759 59703 491775
rect 59669 491683 59703 491699
rect 59827 491759 59861 491775
rect 59827 491683 59861 491699
rect 59945 491759 59979 491775
rect 59945 491683 59979 491699
rect 60103 491759 60137 491775
rect 60103 491683 60137 491699
rect 60221 491759 60255 491775
rect 60221 491683 60255 491699
rect 60379 491759 60413 491775
rect 60379 491683 60413 491699
rect 60497 491759 60531 491775
rect 60497 491683 60531 491699
rect 60655 491759 60689 491775
rect 60655 491683 60689 491699
rect 60773 491759 60807 491775
rect 60773 491683 60807 491699
rect 60931 491759 60965 491775
rect 60931 491683 60965 491699
rect 61049 491759 61083 491775
rect 61049 491683 61083 491699
rect 61207 491759 61241 491775
rect 61207 491683 61241 491699
rect 61325 491759 61359 491775
rect 61325 491683 61359 491699
rect 61483 491759 61517 491775
rect 61483 491683 61517 491699
rect 58904 491649 58982 491650
rect 59730 491649 59808 491650
rect 60006 491649 60084 491650
rect 60278 491649 60356 491652
rect 60556 491649 60634 491650
rect 60834 491649 60912 491652
rect 61110 491649 61188 491652
rect 61386 491649 61464 491654
rect 58887 491615 58903 491649
rect 58971 491615 58987 491649
rect 59163 491615 59179 491649
rect 59247 491615 59263 491649
rect 59439 491615 59455 491649
rect 59523 491615 59539 491649
rect 59715 491615 59731 491649
rect 59799 491615 59815 491649
rect 59991 491615 60007 491649
rect 60075 491615 60091 491649
rect 60267 491615 60283 491649
rect 60351 491615 60367 491649
rect 60543 491615 60559 491649
rect 60627 491615 60643 491649
rect 60819 491615 60835 491649
rect 60903 491615 60919 491649
rect 61095 491615 61111 491649
rect 61179 491615 61195 491649
rect 61371 491615 61387 491649
rect 61455 491615 61471 491649
rect 58904 491514 58982 491615
rect 59178 491514 59256 491615
rect 59454 491514 59532 491615
rect 59730 491514 59808 491615
rect 60006 491608 60084 491615
rect 60278 491514 60356 491615
rect 60556 491514 60634 491615
rect 60834 491514 60912 491615
rect 61110 491514 61188 491615
rect 61386 491514 61464 491615
rect 143336 491780 157833 491838
rect 61617 491557 61651 491573
rect 143335 491740 157833 491780
rect 143335 491553 143422 491740
rect 143620 491553 143718 491740
rect 143896 491553 143994 491740
rect 144170 491553 144268 491740
rect 144448 491553 144546 491740
rect 144720 491553 144818 491740
rect 144998 491553 145096 491740
rect 145276 491553 145374 491740
rect 145554 491553 145652 491740
rect 145828 491553 145926 491740
rect 146104 491553 146202 491740
rect 146389 491553 146484 491740
rect 146658 491553 146756 491740
rect 146934 491553 147032 491740
rect 147206 491553 147304 491740
rect 147484 491553 147582 491740
rect 147756 491553 147854 491740
rect 148034 491553 148132 491740
rect 148310 491553 148408 491740
rect 143335 491530 143353 491553
rect 143337 491519 143353 491530
rect 143421 491519 143437 491553
rect 143613 491519 143629 491553
rect 143697 491529 143718 491553
rect 143697 491519 143713 491529
rect 143889 491519 143905 491553
rect 143973 491531 143994 491553
rect 143973 491519 143989 491531
rect 144165 491519 144181 491553
rect 144249 491527 144268 491553
rect 144249 491519 144265 491527
rect 144441 491519 144457 491553
rect 144525 491527 144546 491553
rect 144525 491519 144541 491527
rect 144717 491519 144733 491553
rect 144801 491529 144818 491553
rect 144801 491519 144817 491529
rect 144993 491519 145009 491553
rect 145077 491527 145096 491553
rect 145077 491519 145093 491527
rect 145269 491519 145285 491553
rect 145353 491527 145374 491553
rect 145353 491519 145369 491527
rect 145545 491519 145561 491553
rect 145629 491531 145652 491553
rect 145629 491519 145645 491531
rect 145821 491519 145837 491553
rect 145905 491527 145926 491553
rect 145905 491519 145921 491527
rect 146097 491519 146113 491553
rect 146181 491531 146202 491553
rect 146181 491519 146197 491531
rect 146373 491519 146389 491553
rect 146457 491530 146484 491553
rect 146457 491519 146473 491530
rect 146649 491519 146665 491553
rect 146733 491533 146756 491553
rect 146733 491519 146749 491533
rect 146925 491519 146941 491553
rect 147009 491523 147032 491553
rect 147009 491519 147025 491523
rect 147201 491519 147217 491553
rect 147285 491527 147304 491553
rect 147285 491519 147301 491527
rect 147477 491519 147493 491553
rect 147561 491527 147582 491553
rect 147561 491519 147577 491527
rect 147753 491519 147769 491553
rect 147837 491519 147854 491553
rect 148029 491519 148045 491553
rect 148113 491527 148132 491553
rect 148113 491519 148129 491527
rect 148305 491519 148321 491553
rect 148389 491527 148408 491553
rect 148580 491553 148678 491740
rect 148866 491553 148964 491740
rect 149138 491553 149236 491740
rect 149418 491553 149516 491740
rect 149692 491553 149790 491740
rect 150244 491553 150342 491740
rect 150520 491553 150618 491740
rect 150796 491553 150894 491740
rect 151072 491553 151170 491740
rect 151348 491553 151446 491740
rect 151624 491553 151722 491740
rect 151902 491553 152000 491740
rect 152178 491553 152276 491740
rect 152450 491553 152548 491740
rect 152728 491553 152826 491740
rect 153004 491553 153102 491740
rect 153282 491553 153380 491740
rect 153556 491553 153654 491740
rect 153832 491553 153930 491740
rect 154110 491553 154208 491740
rect 154386 491553 154484 491740
rect 154662 491553 154760 491740
rect 154938 491553 155036 491740
rect 155214 491553 155312 491740
rect 155488 491553 155586 491740
rect 155768 491553 155866 491740
rect 156044 491553 156142 491740
rect 156316 491553 156414 491740
rect 156592 491553 156690 491740
rect 156862 491553 156960 491740
rect 157154 491553 157252 491740
rect 148389 491519 148405 491527
rect 148580 491525 148597 491553
rect 148581 491519 148597 491525
rect 148665 491519 148681 491553
rect 148857 491519 148873 491553
rect 148941 491523 148964 491553
rect 148941 491519 148957 491523
rect 149133 491519 149149 491553
rect 149217 491523 149236 491553
rect 149217 491519 149233 491523
rect 149409 491519 149425 491553
rect 149493 491523 149516 491553
rect 149493 491519 149509 491523
rect 149685 491519 149701 491553
rect 149769 491523 149790 491553
rect 149769 491519 149785 491523
rect 149961 491519 149977 491553
rect 150045 491519 150061 491553
rect 150237 491519 150253 491553
rect 150321 491523 150342 491553
rect 150321 491519 150337 491523
rect 150513 491519 150529 491553
rect 150597 491525 150618 491553
rect 150597 491519 150613 491525
rect 150789 491519 150805 491553
rect 150873 491525 150894 491553
rect 150873 491519 150889 491525
rect 151065 491519 151081 491553
rect 151149 491527 151170 491553
rect 151149 491519 151165 491527
rect 151341 491519 151357 491553
rect 151425 491525 151446 491553
rect 151425 491519 151441 491525
rect 151617 491519 151633 491553
rect 151701 491525 151722 491553
rect 151701 491519 151717 491525
rect 151893 491519 151909 491553
rect 151977 491525 152000 491553
rect 151977 491519 151993 491525
rect 152169 491519 152185 491553
rect 152253 491525 152276 491553
rect 152253 491519 152269 491525
rect 152445 491519 152461 491553
rect 152529 491523 152548 491553
rect 152529 491519 152545 491523
rect 152721 491519 152737 491553
rect 152805 491523 152826 491553
rect 152805 491519 152821 491523
rect 152997 491519 153013 491553
rect 153081 491527 153102 491553
rect 153081 491519 153097 491527
rect 153273 491519 153289 491553
rect 153357 491529 153380 491553
rect 153357 491519 153373 491529
rect 153549 491519 153565 491553
rect 153633 491525 153654 491553
rect 153633 491519 153649 491525
rect 153825 491519 153841 491553
rect 153909 491529 153930 491553
rect 153909 491519 153925 491529
rect 154101 491519 154117 491553
rect 154185 491529 154208 491553
rect 154185 491519 154201 491529
rect 154377 491519 154393 491553
rect 154461 491531 154484 491553
rect 154461 491519 154477 491531
rect 154653 491519 154669 491553
rect 154737 491527 154760 491553
rect 154737 491519 154753 491527
rect 154929 491519 154945 491553
rect 155013 491529 155036 491553
rect 155013 491519 155029 491529
rect 155205 491519 155221 491553
rect 155289 491529 155312 491553
rect 155289 491519 155305 491529
rect 155481 491519 155497 491553
rect 155565 491531 155586 491553
rect 155565 491519 155581 491531
rect 155757 491519 155773 491553
rect 155841 491531 155866 491553
rect 155841 491519 155857 491531
rect 156033 491519 156049 491553
rect 156117 491531 156142 491553
rect 156117 491519 156133 491531
rect 156309 491519 156325 491553
rect 156393 491531 156414 491553
rect 156393 491519 156409 491531
rect 156585 491519 156601 491553
rect 156669 491521 156690 491553
rect 156669 491519 156685 491521
rect 156861 491519 156877 491553
rect 156945 491519 156961 491553
rect 157137 491519 157153 491553
rect 157221 491521 157252 491553
rect 157383 491595 157417 491611
rect 157221 491519 157237 491521
rect 58580 491472 61466 491514
rect 59544 491334 59660 491472
rect 143291 491469 143325 491485
rect 143291 491393 143325 491409
rect 143449 491469 143483 491485
rect 143449 491393 143483 491409
rect 143567 491469 143601 491485
rect 143567 491393 143601 491409
rect 143725 491469 143759 491485
rect 143725 491393 143759 491409
rect 143843 491469 143877 491485
rect 143843 491393 143877 491409
rect 144001 491469 144035 491485
rect 144001 491393 144035 491409
rect 144119 491469 144153 491485
rect 144119 491393 144153 491409
rect 144277 491469 144311 491485
rect 144277 491393 144311 491409
rect 144395 491469 144429 491485
rect 144395 491393 144429 491409
rect 144553 491469 144587 491485
rect 144553 491393 144587 491409
rect 144671 491469 144705 491485
rect 144671 491393 144705 491409
rect 144829 491469 144863 491485
rect 144829 491393 144863 491409
rect 144947 491469 144981 491485
rect 144947 491393 144981 491409
rect 145105 491469 145139 491485
rect 145105 491393 145139 491409
rect 145223 491469 145257 491485
rect 145223 491393 145257 491409
rect 145381 491469 145415 491485
rect 145381 491393 145415 491409
rect 145499 491469 145533 491485
rect 145499 491393 145533 491409
rect 145657 491469 145691 491485
rect 145657 491393 145691 491409
rect 145775 491469 145809 491485
rect 145775 491393 145809 491409
rect 145933 491469 145967 491485
rect 145933 491393 145967 491409
rect 146051 491469 146085 491485
rect 146051 491393 146085 491409
rect 146209 491469 146243 491485
rect 146209 491393 146243 491409
rect 146327 491469 146361 491485
rect 146327 491393 146361 491409
rect 146485 491469 146519 491485
rect 146485 491393 146519 491409
rect 146603 491469 146637 491485
rect 146603 491393 146637 491409
rect 146761 491469 146795 491485
rect 146761 491393 146795 491409
rect 146879 491469 146913 491485
rect 146879 491393 146913 491409
rect 147037 491469 147071 491485
rect 147037 491393 147071 491409
rect 147155 491469 147189 491485
rect 147155 491393 147189 491409
rect 147313 491469 147347 491485
rect 147313 491393 147347 491409
rect 147431 491469 147465 491485
rect 147431 491393 147465 491409
rect 147589 491469 147623 491485
rect 147589 491393 147623 491409
rect 147707 491469 147741 491485
rect 147707 491393 147741 491409
rect 147865 491469 147899 491485
rect 147865 491393 147899 491409
rect 147983 491469 148017 491485
rect 147983 491393 148017 491409
rect 148141 491469 148175 491485
rect 148141 491393 148175 491409
rect 148259 491469 148293 491485
rect 148259 491393 148293 491409
rect 148417 491469 148451 491485
rect 148417 491393 148451 491409
rect 148535 491469 148569 491485
rect 148535 491393 148569 491409
rect 148693 491469 148727 491485
rect 148693 491393 148727 491409
rect 148811 491469 148845 491485
rect 148811 491393 148845 491409
rect 148969 491469 149003 491485
rect 148969 491393 149003 491409
rect 149087 491469 149121 491485
rect 149087 491393 149121 491409
rect 149245 491469 149279 491485
rect 149245 491393 149279 491409
rect 149363 491469 149397 491485
rect 149363 491393 149397 491409
rect 149521 491469 149555 491485
rect 149521 491393 149555 491409
rect 149639 491469 149673 491485
rect 149639 491393 149673 491409
rect 149797 491469 149831 491485
rect 149797 491393 149831 491409
rect 149915 491469 149949 491485
rect 149915 491393 149949 491409
rect 150073 491469 150107 491485
rect 150073 491393 150107 491409
rect 150191 491469 150225 491485
rect 150191 491393 150225 491409
rect 150349 491469 150383 491485
rect 150349 491393 150383 491409
rect 150467 491469 150501 491485
rect 150467 491393 150501 491409
rect 150625 491469 150659 491485
rect 150625 491393 150659 491409
rect 150743 491469 150777 491485
rect 150743 491393 150777 491409
rect 150901 491469 150935 491485
rect 150901 491393 150935 491409
rect 151019 491469 151053 491485
rect 151019 491393 151053 491409
rect 151177 491469 151211 491485
rect 151177 491393 151211 491409
rect 151295 491469 151329 491485
rect 151295 491393 151329 491409
rect 151453 491469 151487 491485
rect 151453 491393 151487 491409
rect 151571 491469 151605 491485
rect 151571 491393 151605 491409
rect 151729 491469 151763 491485
rect 151729 491393 151763 491409
rect 151847 491469 151881 491485
rect 151847 491393 151881 491409
rect 152005 491469 152039 491485
rect 152005 491393 152039 491409
rect 152123 491469 152157 491485
rect 152123 491393 152157 491409
rect 152281 491469 152315 491485
rect 152281 491393 152315 491409
rect 152399 491469 152433 491485
rect 152399 491393 152433 491409
rect 152557 491469 152591 491485
rect 152557 491393 152591 491409
rect 152675 491469 152709 491485
rect 152675 491393 152709 491409
rect 152833 491469 152867 491485
rect 152833 491393 152867 491409
rect 152951 491469 152985 491485
rect 152951 491393 152985 491409
rect 153109 491469 153143 491485
rect 153109 491393 153143 491409
rect 153227 491469 153261 491485
rect 153227 491393 153261 491409
rect 153385 491469 153419 491485
rect 153385 491393 153419 491409
rect 153503 491469 153537 491485
rect 153503 491393 153537 491409
rect 153661 491469 153695 491485
rect 153661 491393 153695 491409
rect 153779 491469 153813 491485
rect 153779 491393 153813 491409
rect 153937 491469 153971 491485
rect 153937 491393 153971 491409
rect 154055 491469 154089 491485
rect 154055 491393 154089 491409
rect 154213 491469 154247 491485
rect 154213 491393 154247 491409
rect 154331 491469 154365 491485
rect 154331 491393 154365 491409
rect 154489 491469 154523 491485
rect 154489 491393 154523 491409
rect 154607 491469 154641 491485
rect 154607 491393 154641 491409
rect 154765 491469 154799 491485
rect 154765 491393 154799 491409
rect 154883 491469 154917 491485
rect 154883 491393 154917 491409
rect 155041 491469 155075 491485
rect 155041 491393 155075 491409
rect 155159 491469 155193 491485
rect 155159 491393 155193 491409
rect 155317 491469 155351 491485
rect 155317 491393 155351 491409
rect 155435 491469 155469 491485
rect 155435 491393 155469 491409
rect 155593 491469 155627 491485
rect 155593 491393 155627 491409
rect 155711 491469 155745 491485
rect 155711 491393 155745 491409
rect 155869 491469 155903 491485
rect 155869 491393 155903 491409
rect 155987 491469 156021 491485
rect 155987 491393 156021 491409
rect 156145 491469 156179 491485
rect 156145 491393 156179 491409
rect 156263 491469 156297 491485
rect 156263 491393 156297 491409
rect 156421 491469 156455 491485
rect 156421 491393 156455 491409
rect 156539 491469 156573 491485
rect 156539 491393 156573 491409
rect 156697 491469 156731 491485
rect 156697 491393 156731 491409
rect 156815 491469 156849 491485
rect 156815 491393 156849 491409
rect 156973 491469 157007 491485
rect 156973 491393 157007 491409
rect 157091 491469 157125 491485
rect 157091 491393 157125 491409
rect 157249 491469 157283 491485
rect 157249 491393 157283 491409
rect 59544 491290 59566 491334
rect 59638 491290 59660 491334
rect 143337 491325 143353 491359
rect 143421 491356 143437 491359
rect 143421 491325 143445 491356
rect 143613 491325 143629 491359
rect 143697 491325 143713 491359
rect 143889 491355 143905 491359
rect 143886 491325 143905 491355
rect 143973 491325 143989 491359
rect 144165 491351 144181 491359
rect 144162 491325 144181 491351
rect 144249 491325 144265 491359
rect 144441 491345 144457 491359
rect 144440 491325 144457 491345
rect 144525 491325 144541 491359
rect 144717 491341 144733 491359
rect 144716 491325 144733 491341
rect 144801 491325 144817 491359
rect 144993 491343 145009 491359
rect 144990 491325 145009 491343
rect 145077 491325 145093 491359
rect 145269 491341 145285 491359
rect 145268 491325 145285 491341
rect 145353 491325 145369 491359
rect 145545 491325 145561 491359
rect 145629 491325 145645 491359
rect 145821 491341 145837 491359
rect 145820 491325 145837 491341
rect 145905 491325 145921 491359
rect 146097 491325 146113 491359
rect 146181 491325 146197 491359
rect 146373 491351 146389 491359
rect 146370 491335 146389 491351
rect 146369 491325 146389 491335
rect 146457 491325 146473 491359
rect 146649 491351 146665 491359
rect 146646 491325 146665 491351
rect 146733 491325 146749 491359
rect 146925 491325 146941 491359
rect 147009 491325 147025 491359
rect 147201 491345 147217 491359
rect 147194 491325 147217 491345
rect 147285 491325 147301 491359
rect 147477 491325 147493 491359
rect 147561 491325 147577 491359
rect 147753 491345 147769 491359
rect 147752 491325 147769 491345
rect 147837 491325 147853 491359
rect 148029 491341 148045 491359
rect 148028 491325 148045 491341
rect 148113 491325 148129 491359
rect 148305 491349 148321 491359
rect 148302 491325 148321 491349
rect 148389 491325 148405 491359
rect 148581 491341 148597 491359
rect 148580 491325 148597 491341
rect 148665 491325 148681 491359
rect 148857 491343 148873 491359
rect 148850 491325 148873 491343
rect 148941 491325 148957 491359
rect 149133 491349 149149 491359
rect 149126 491325 149149 491349
rect 149217 491325 149233 491359
rect 149409 491355 149425 491359
rect 149408 491325 149425 491355
rect 149493 491325 149509 491359
rect 149685 491351 149701 491359
rect 149684 491325 149701 491351
rect 149769 491325 149785 491359
rect 149961 491351 149977 491359
rect 149958 491325 149977 491351
rect 150045 491325 150061 491359
rect 150237 491351 150253 491359
rect 150230 491325 150253 491351
rect 150321 491325 150337 491359
rect 150513 491351 150529 491359
rect 150512 491325 150529 491351
rect 150597 491325 150613 491359
rect 150789 491325 150805 491359
rect 150873 491325 150889 491359
rect 151065 491345 151081 491359
rect 151064 491325 151081 491345
rect 151149 491325 151165 491359
rect 151341 491325 151357 491359
rect 151425 491325 151441 491359
rect 151617 491325 151633 491359
rect 151701 491325 151717 491359
rect 151893 491337 151909 491359
rect 151886 491325 151909 491337
rect 151977 491325 151993 491359
rect 152169 491333 152185 491359
rect 152168 491325 152185 491333
rect 152253 491325 152269 491359
rect 152445 491325 152461 491359
rect 152529 491325 152545 491359
rect 152721 491333 152737 491359
rect 152720 491325 152737 491333
rect 152805 491325 152821 491359
rect 152997 491333 153013 491359
rect 152996 491325 153013 491333
rect 153081 491325 153097 491359
rect 153273 491349 153289 491359
rect 153266 491325 153289 491349
rect 153357 491325 153373 491359
rect 153549 491341 153565 491359
rect 153544 491325 153565 491341
rect 153633 491325 153649 491359
rect 153825 491325 153841 491359
rect 153909 491325 153925 491359
rect 154101 491325 154117 491359
rect 154185 491341 154201 491359
rect 154377 491345 154393 491359
rect 154185 491325 154206 491341
rect 59544 491264 59660 491290
rect 59602 491258 59660 491264
rect 143343 491116 143445 491325
rect 143614 491116 143712 491325
rect 143886 491116 143984 491325
rect 144162 491116 144260 491325
rect 144440 491116 144538 491325
rect 144716 491116 144814 491325
rect 144990 491116 145088 491325
rect 145268 491116 145366 491325
rect 145546 491116 145644 491325
rect 145820 491116 145918 491325
rect 146098 491116 146196 491325
rect 146369 491116 146469 491325
rect 146646 491116 146744 491325
rect 146926 491116 147024 491325
rect 147194 491116 147292 491325
rect 147478 491116 147576 491325
rect 147752 491116 147850 491325
rect 148028 491116 148126 491325
rect 148302 491116 148400 491325
rect 148580 491116 148678 491325
rect 148850 491116 148948 491325
rect 149126 491116 149224 491325
rect 149408 491116 149506 491325
rect 149684 491116 149782 491325
rect 149958 491310 150056 491325
rect 150230 491116 150328 491325
rect 150512 491116 150610 491325
rect 150790 491116 150888 491325
rect 151064 491116 151162 491325
rect 151342 491116 151440 491325
rect 151618 491116 151716 491325
rect 151886 491116 151984 491325
rect 152168 491116 152266 491325
rect 152446 491116 152544 491325
rect 152720 491116 152818 491325
rect 152996 491116 153094 491325
rect 153266 491116 153364 491325
rect 153544 491116 153642 491325
rect 153826 491116 153924 491325
rect 154108 491116 154206 491325
rect 154376 491325 154393 491345
rect 154461 491325 154477 491359
rect 154653 491345 154669 491359
rect 154652 491325 154669 491345
rect 154737 491325 154753 491359
rect 154929 491345 154945 491359
rect 154922 491325 154945 491345
rect 155013 491325 155029 491359
rect 155205 491351 155221 491359
rect 155200 491325 155221 491351
rect 155289 491325 155305 491359
rect 155481 491325 155497 491359
rect 155565 491325 155581 491359
rect 155757 491325 155773 491359
rect 155841 491351 155857 491359
rect 155841 491325 155860 491351
rect 156033 491349 156049 491359
rect 154376 491116 154474 491325
rect 154652 491116 154750 491325
rect 154922 491116 155020 491325
rect 155200 491116 155298 491325
rect 155482 491116 155580 491325
rect 155762 491116 155860 491325
rect 156028 491325 156049 491349
rect 156117 491325 156133 491359
rect 156309 491343 156325 491359
rect 156304 491325 156325 491343
rect 156393 491325 156409 491359
rect 156585 491349 156601 491359
rect 156584 491325 156601 491349
rect 156669 491325 156685 491359
rect 156861 491325 156877 491359
rect 156945 491349 156961 491359
rect 156945 491325 156966 491349
rect 157137 491325 157153 491359
rect 157221 491353 157237 491359
rect 157221 491325 157244 491353
rect 156028 491116 156126 491325
rect 156304 491116 156402 491325
rect 156584 491116 156682 491325
rect 156868 491116 156966 491325
rect 157146 491116 157244 491325
rect 157383 491267 157417 491283
rect 157735 491116 157833 491740
rect 323888 491686 323968 492003
rect 324154 491793 324252 492003
rect 324426 491793 324524 492003
rect 324702 491793 324800 492003
rect 324980 491793 325078 492003
rect 325256 491793 325354 492003
rect 325530 491793 325628 492003
rect 325808 491793 325906 492003
rect 326086 491793 326184 492003
rect 326360 491793 326458 492003
rect 326638 491793 326736 492003
rect 326910 491793 327008 492003
rect 327186 491793 327284 492003
rect 327466 491793 327564 492003
rect 327734 491793 327832 492003
rect 328018 491793 328116 492003
rect 328292 491793 328390 492003
rect 328568 491793 328666 492003
rect 328842 491793 328940 492003
rect 329120 491793 329218 492003
rect 329390 491793 329488 492003
rect 329666 491793 329764 492003
rect 329948 491793 330046 492003
rect 330224 491793 330322 492003
rect 330498 491793 330596 492003
rect 330770 491793 330868 492003
rect 331052 491793 331150 492003
rect 331330 491793 331428 492003
rect 331604 491793 331702 492003
rect 331882 491793 331980 492003
rect 332158 491793 332256 492003
rect 332426 491793 332524 492003
rect 332708 491793 332806 492003
rect 332986 491793 333084 492003
rect 333260 491793 333358 492003
rect 333536 491793 333634 492003
rect 333806 491793 333904 492003
rect 334084 491793 334182 492003
rect 334366 491793 334464 492003
rect 334648 491793 334746 492003
rect 334916 492003 334933 492022
rect 335001 492003 335017 492037
rect 335193 492022 335209 492037
rect 335192 492003 335209 492022
rect 335277 492003 335293 492037
rect 335469 492022 335485 492037
rect 335462 492003 335485 492022
rect 335553 492003 335569 492037
rect 335745 492028 335761 492037
rect 335740 492003 335761 492028
rect 335829 492003 335845 492037
rect 336021 492003 336037 492037
rect 336105 492003 336121 492037
rect 336297 492003 336313 492037
rect 336381 492028 336397 492037
rect 336381 492003 336400 492028
rect 336573 492026 336589 492037
rect 334916 491793 335014 492003
rect 335192 491793 335290 492003
rect 335462 491793 335560 492003
rect 335740 491793 335838 492003
rect 336022 491793 336120 492003
rect 336302 491793 336400 492003
rect 336568 492003 336589 492026
rect 336657 492003 336673 492037
rect 336849 492020 336865 492037
rect 336844 492003 336865 492020
rect 336933 492003 336949 492037
rect 337125 492026 337141 492037
rect 337124 492003 337141 492026
rect 337209 492003 337225 492037
rect 337401 492003 337417 492037
rect 337485 492026 337501 492037
rect 337485 492003 337506 492026
rect 337677 492003 337693 492037
rect 337761 492030 337777 492037
rect 337761 492003 337784 492030
rect 336568 491793 336666 492003
rect 336844 491793 336942 492003
rect 337124 491793 337222 492003
rect 337408 491793 337506 492003
rect 337686 491793 337784 492003
rect 337923 491945 337957 491961
rect 338275 491793 338373 492417
rect 324154 491762 338373 491793
rect 324154 491706 327886 491762
rect 327964 491706 338373 491762
rect 324154 491695 338373 491706
rect 508580 491988 511459 491999
rect 508580 491957 511460 491988
rect 323888 491644 323904 491686
rect 323958 491644 323968 491686
rect 323888 491624 323968 491644
rect 418707 491582 420075 491618
rect 418707 491246 418743 491582
rect 418907 491515 418977 491582
rect 419175 491515 419245 491582
rect 419723 491515 419793 491582
rect 420005 491515 420075 491582
rect 420236 491557 420270 491573
rect 418886 491481 418902 491515
rect 418970 491481 418986 491515
rect 419162 491481 419178 491515
rect 419246 491481 419262 491515
rect 419438 491481 419454 491515
rect 419522 491481 419538 491515
rect 419714 491481 419730 491515
rect 419798 491481 419814 491515
rect 419990 491481 420006 491515
rect 420074 491481 420090 491515
rect 418907 491476 418977 491481
rect 419175 491476 419245 491481
rect 419723 491474 419793 491481
rect 420005 491476 420075 491481
rect 418840 491431 418874 491447
rect 418840 491355 418874 491371
rect 418998 491431 419032 491447
rect 418998 491355 419032 491371
rect 419116 491431 419150 491447
rect 419116 491355 419150 491371
rect 419274 491431 419308 491447
rect 419274 491355 419308 491371
rect 419392 491431 419426 491447
rect 419392 491355 419426 491371
rect 419550 491431 419584 491447
rect 419550 491355 419584 491371
rect 419668 491431 419702 491447
rect 419668 491355 419702 491371
rect 419826 491431 419860 491447
rect 419826 491355 419860 491371
rect 419944 491431 419978 491447
rect 419944 491355 419978 491371
rect 420102 491431 420136 491447
rect 420102 491355 420136 491371
rect 419721 491321 419817 491322
rect 418886 491287 418902 491321
rect 418970 491287 418986 491321
rect 419162 491287 419178 491321
rect 419246 491287 419262 491321
rect 419438 491287 419454 491321
rect 419522 491287 419538 491321
rect 419714 491287 419730 491321
rect 419798 491287 419817 491321
rect 419990 491287 420006 491321
rect 420074 491287 420090 491321
rect 419165 491246 419259 491287
rect 419721 491250 419817 491287
rect 420011 491260 420075 491287
rect 420011 491250 420073 491260
rect 419719 491246 420073 491250
rect 418707 491244 420073 491246
rect 232693 491184 247190 491242
rect 418707 491210 418923 491244
rect 418961 491210 420073 491244
rect 508580 491514 508622 491957
rect 508900 491952 511460 491957
rect 508900 491843 508978 491952
rect 509176 491843 509254 491952
rect 509454 491843 509532 491952
rect 509726 491843 509804 491952
rect 510008 491843 510086 491850
rect 510280 491843 510358 491952
rect 510556 491843 510634 491952
rect 510830 491843 510908 491952
rect 511108 491843 511186 491952
rect 511382 491843 511460 491952
rect 511617 491885 511651 491901
rect 508887 491809 508903 491843
rect 508971 491809 508987 491843
rect 509163 491809 509179 491843
rect 509247 491809 509263 491843
rect 509439 491809 509455 491843
rect 509523 491809 509539 491843
rect 509715 491809 509731 491843
rect 509799 491809 509815 491843
rect 509991 491809 510007 491843
rect 510075 491809 510091 491843
rect 510267 491809 510283 491843
rect 510351 491809 510367 491843
rect 510543 491809 510559 491843
rect 510627 491809 510643 491843
rect 510819 491809 510835 491843
rect 510903 491809 510919 491843
rect 511095 491809 511111 491843
rect 511179 491809 511195 491843
rect 511371 491809 511387 491843
rect 511455 491809 511471 491843
rect 508900 491808 508978 491809
rect 509176 491806 509254 491809
rect 509454 491808 509532 491809
rect 509726 491808 509804 491809
rect 510008 491808 510086 491809
rect 510280 491808 510358 491809
rect 510556 491806 510634 491809
rect 510830 491806 510908 491809
rect 511108 491808 511186 491809
rect 511382 491806 511460 491809
rect 508841 491759 508875 491775
rect 508841 491683 508875 491699
rect 508999 491759 509033 491775
rect 508999 491683 509033 491699
rect 509117 491759 509151 491775
rect 509117 491683 509151 491699
rect 509275 491759 509309 491775
rect 509275 491683 509309 491699
rect 509393 491759 509427 491775
rect 509393 491683 509427 491699
rect 509551 491759 509585 491775
rect 509551 491683 509585 491699
rect 509669 491759 509703 491775
rect 509669 491683 509703 491699
rect 509827 491759 509861 491775
rect 509827 491683 509861 491699
rect 509945 491759 509979 491775
rect 509945 491683 509979 491699
rect 510103 491759 510137 491775
rect 510103 491683 510137 491699
rect 510221 491759 510255 491775
rect 510221 491683 510255 491699
rect 510379 491759 510413 491775
rect 510379 491683 510413 491699
rect 510497 491759 510531 491775
rect 510497 491683 510531 491699
rect 510655 491759 510689 491775
rect 510655 491683 510689 491699
rect 510773 491759 510807 491775
rect 510773 491683 510807 491699
rect 510931 491759 510965 491775
rect 510931 491683 510965 491699
rect 511049 491759 511083 491775
rect 511049 491683 511083 491699
rect 511207 491759 511241 491775
rect 511207 491683 511241 491699
rect 511325 491759 511359 491775
rect 511325 491683 511359 491699
rect 511483 491759 511517 491775
rect 511483 491683 511517 491699
rect 508904 491649 508982 491650
rect 509730 491649 509808 491650
rect 510006 491649 510084 491650
rect 510278 491649 510356 491652
rect 510556 491649 510634 491650
rect 510834 491649 510912 491652
rect 511110 491649 511188 491652
rect 511386 491649 511464 491654
rect 508887 491615 508903 491649
rect 508971 491615 508987 491649
rect 509163 491615 509179 491649
rect 509247 491615 509263 491649
rect 509439 491615 509455 491649
rect 509523 491615 509539 491649
rect 509715 491615 509731 491649
rect 509799 491615 509815 491649
rect 509991 491615 510007 491649
rect 510075 491615 510091 491649
rect 510267 491615 510283 491649
rect 510351 491615 510367 491649
rect 510543 491615 510559 491649
rect 510627 491615 510643 491649
rect 510819 491615 510835 491649
rect 510903 491615 510919 491649
rect 511095 491615 511111 491649
rect 511179 491615 511195 491649
rect 511371 491615 511387 491649
rect 511455 491615 511471 491649
rect 508904 491514 508982 491615
rect 509178 491514 509256 491615
rect 509454 491514 509532 491615
rect 509730 491514 509808 491615
rect 510006 491608 510084 491615
rect 510278 491514 510356 491615
rect 510556 491514 510634 491615
rect 510834 491514 510912 491615
rect 511110 491514 511188 491615
rect 511386 491514 511464 491615
rect 511617 491557 511651 491573
rect 508580 491472 511466 491514
rect 509544 491334 509660 491472
rect 509544 491290 509566 491334
rect 509638 491290 509660 491334
rect 509544 491264 509660 491290
rect 509602 491258 509660 491264
rect 420236 491229 420270 491245
rect 419719 491208 420073 491210
rect 143340 491085 157833 491116
rect 143340 491029 147346 491085
rect 147424 491029 157833 491085
rect 143340 491018 157833 491029
rect 232692 491144 247190 491184
rect 232692 490957 232779 491144
rect 232977 490957 233075 491144
rect 233253 490957 233351 491144
rect 233527 490957 233625 491144
rect 233805 490957 233903 491144
rect 234077 490957 234175 491144
rect 234355 490957 234453 491144
rect 234633 490957 234731 491144
rect 234911 490957 235009 491144
rect 235185 490957 235283 491144
rect 235461 490957 235559 491144
rect 235746 490957 235841 491144
rect 236015 490957 236113 491144
rect 236291 490957 236389 491144
rect 236563 490957 236661 491144
rect 236841 490957 236939 491144
rect 237113 490957 237211 491144
rect 237391 490957 237489 491144
rect 237667 490957 237765 491144
rect 232692 490934 232710 490957
rect 232694 490923 232710 490934
rect 232778 490923 232794 490957
rect 232970 490923 232986 490957
rect 233054 490933 233075 490957
rect 233054 490923 233070 490933
rect 233246 490923 233262 490957
rect 233330 490935 233351 490957
rect 233330 490923 233346 490935
rect 233522 490923 233538 490957
rect 233606 490931 233625 490957
rect 233606 490923 233622 490931
rect 233798 490923 233814 490957
rect 233882 490931 233903 490957
rect 233882 490923 233898 490931
rect 234074 490923 234090 490957
rect 234158 490933 234175 490957
rect 234158 490923 234174 490933
rect 234350 490923 234366 490957
rect 234434 490931 234453 490957
rect 234434 490923 234450 490931
rect 234626 490923 234642 490957
rect 234710 490931 234731 490957
rect 234710 490923 234726 490931
rect 234902 490923 234918 490957
rect 234986 490935 235009 490957
rect 234986 490923 235002 490935
rect 235178 490923 235194 490957
rect 235262 490931 235283 490957
rect 235262 490923 235278 490931
rect 235454 490923 235470 490957
rect 235538 490935 235559 490957
rect 235538 490923 235554 490935
rect 235730 490923 235746 490957
rect 235814 490934 235841 490957
rect 235814 490923 235830 490934
rect 236006 490923 236022 490957
rect 236090 490937 236113 490957
rect 236090 490923 236106 490937
rect 236282 490923 236298 490957
rect 236366 490927 236389 490957
rect 236366 490923 236382 490927
rect 236558 490923 236574 490957
rect 236642 490931 236661 490957
rect 236642 490923 236658 490931
rect 236834 490923 236850 490957
rect 236918 490931 236939 490957
rect 236918 490923 236934 490931
rect 237110 490923 237126 490957
rect 237194 490923 237211 490957
rect 237386 490923 237402 490957
rect 237470 490931 237489 490957
rect 237470 490923 237486 490931
rect 237662 490923 237678 490957
rect 237746 490931 237765 490957
rect 237937 490957 238035 491144
rect 238223 490957 238321 491144
rect 238495 490957 238593 491144
rect 238775 490957 238873 491144
rect 239049 490957 239147 491144
rect 239601 490957 239699 491144
rect 239877 490957 239975 491144
rect 240153 490957 240251 491144
rect 240429 490957 240527 491144
rect 240705 490957 240803 491144
rect 240981 490957 241079 491144
rect 241259 490957 241357 491144
rect 241535 490957 241633 491144
rect 241807 490957 241905 491144
rect 242085 490957 242183 491144
rect 242361 490957 242459 491144
rect 242639 490957 242737 491144
rect 242913 490957 243011 491144
rect 243189 490957 243287 491144
rect 243467 490957 243565 491144
rect 243743 490957 243841 491144
rect 244019 490957 244117 491144
rect 244295 490957 244393 491144
rect 244571 490957 244669 491144
rect 244845 490957 244943 491144
rect 245125 490957 245223 491144
rect 245401 490957 245499 491144
rect 245673 490957 245771 491144
rect 245949 490957 246047 491144
rect 246219 490957 246317 491144
rect 246511 490957 246609 491144
rect 237746 490923 237762 490931
rect 237937 490929 237954 490957
rect 237938 490923 237954 490929
rect 238022 490923 238038 490957
rect 238214 490923 238230 490957
rect 238298 490927 238321 490957
rect 238298 490923 238314 490927
rect 238490 490923 238506 490957
rect 238574 490927 238593 490957
rect 238574 490923 238590 490927
rect 238766 490923 238782 490957
rect 238850 490927 238873 490957
rect 238850 490923 238866 490927
rect 239042 490923 239058 490957
rect 239126 490927 239147 490957
rect 239126 490923 239142 490927
rect 239318 490923 239334 490957
rect 239402 490923 239418 490957
rect 239594 490923 239610 490957
rect 239678 490927 239699 490957
rect 239678 490923 239694 490927
rect 239870 490923 239886 490957
rect 239954 490929 239975 490957
rect 239954 490923 239970 490929
rect 240146 490923 240162 490957
rect 240230 490929 240251 490957
rect 240230 490923 240246 490929
rect 240422 490923 240438 490957
rect 240506 490931 240527 490957
rect 240506 490923 240522 490931
rect 240698 490923 240714 490957
rect 240782 490929 240803 490957
rect 240782 490923 240798 490929
rect 240974 490923 240990 490957
rect 241058 490929 241079 490957
rect 241058 490923 241074 490929
rect 241250 490923 241266 490957
rect 241334 490929 241357 490957
rect 241334 490923 241350 490929
rect 241526 490923 241542 490957
rect 241610 490929 241633 490957
rect 241610 490923 241626 490929
rect 241802 490923 241818 490957
rect 241886 490927 241905 490957
rect 241886 490923 241902 490927
rect 242078 490923 242094 490957
rect 242162 490927 242183 490957
rect 242162 490923 242178 490927
rect 242354 490923 242370 490957
rect 242438 490931 242459 490957
rect 242438 490923 242454 490931
rect 242630 490923 242646 490957
rect 242714 490933 242737 490957
rect 242714 490923 242730 490933
rect 242906 490923 242922 490957
rect 242990 490929 243011 490957
rect 242990 490923 243006 490929
rect 243182 490923 243198 490957
rect 243266 490933 243287 490957
rect 243266 490923 243282 490933
rect 243458 490923 243474 490957
rect 243542 490933 243565 490957
rect 243542 490923 243558 490933
rect 243734 490923 243750 490957
rect 243818 490935 243841 490957
rect 243818 490923 243834 490935
rect 244010 490923 244026 490957
rect 244094 490931 244117 490957
rect 244094 490923 244110 490931
rect 244286 490923 244302 490957
rect 244370 490933 244393 490957
rect 244370 490923 244386 490933
rect 244562 490923 244578 490957
rect 244646 490933 244669 490957
rect 244646 490923 244662 490933
rect 244838 490923 244854 490957
rect 244922 490935 244943 490957
rect 244922 490923 244938 490935
rect 245114 490923 245130 490957
rect 245198 490935 245223 490957
rect 245198 490923 245214 490935
rect 245390 490923 245406 490957
rect 245474 490935 245499 490957
rect 245474 490923 245490 490935
rect 245666 490923 245682 490957
rect 245750 490935 245771 490957
rect 245750 490923 245766 490935
rect 245942 490923 245958 490957
rect 246026 490925 246047 490957
rect 246026 490923 246042 490925
rect 246218 490923 246234 490957
rect 246302 490923 246318 490957
rect 246494 490923 246510 490957
rect 246578 490925 246609 490957
rect 246740 490999 246774 491015
rect 246578 490923 246594 490925
rect 232648 490873 232682 490889
rect 232648 490797 232682 490813
rect 232806 490873 232840 490889
rect 232806 490797 232840 490813
rect 232924 490873 232958 490889
rect 232924 490797 232958 490813
rect 233082 490873 233116 490889
rect 233082 490797 233116 490813
rect 233200 490873 233234 490889
rect 233200 490797 233234 490813
rect 233358 490873 233392 490889
rect 233358 490797 233392 490813
rect 233476 490873 233510 490889
rect 233476 490797 233510 490813
rect 233634 490873 233668 490889
rect 233634 490797 233668 490813
rect 233752 490873 233786 490889
rect 233752 490797 233786 490813
rect 233910 490873 233944 490889
rect 233910 490797 233944 490813
rect 234028 490873 234062 490889
rect 234028 490797 234062 490813
rect 234186 490873 234220 490889
rect 234186 490797 234220 490813
rect 234304 490873 234338 490889
rect 234304 490797 234338 490813
rect 234462 490873 234496 490889
rect 234462 490797 234496 490813
rect 234580 490873 234614 490889
rect 234580 490797 234614 490813
rect 234738 490873 234772 490889
rect 234738 490797 234772 490813
rect 234856 490873 234890 490889
rect 234856 490797 234890 490813
rect 235014 490873 235048 490889
rect 235014 490797 235048 490813
rect 235132 490873 235166 490889
rect 235132 490797 235166 490813
rect 235290 490873 235324 490889
rect 235290 490797 235324 490813
rect 235408 490873 235442 490889
rect 235408 490797 235442 490813
rect 235566 490873 235600 490889
rect 235566 490797 235600 490813
rect 235684 490873 235718 490889
rect 235684 490797 235718 490813
rect 235842 490873 235876 490889
rect 235842 490797 235876 490813
rect 235960 490873 235994 490889
rect 235960 490797 235994 490813
rect 236118 490873 236152 490889
rect 236118 490797 236152 490813
rect 236236 490873 236270 490889
rect 236236 490797 236270 490813
rect 236394 490873 236428 490889
rect 236394 490797 236428 490813
rect 236512 490873 236546 490889
rect 236512 490797 236546 490813
rect 236670 490873 236704 490889
rect 236670 490797 236704 490813
rect 236788 490873 236822 490889
rect 236788 490797 236822 490813
rect 236946 490873 236980 490889
rect 236946 490797 236980 490813
rect 237064 490873 237098 490889
rect 237064 490797 237098 490813
rect 237222 490873 237256 490889
rect 237222 490797 237256 490813
rect 237340 490873 237374 490889
rect 237340 490797 237374 490813
rect 237498 490873 237532 490889
rect 237498 490797 237532 490813
rect 237616 490873 237650 490889
rect 237616 490797 237650 490813
rect 237774 490873 237808 490889
rect 237774 490797 237808 490813
rect 237892 490873 237926 490889
rect 237892 490797 237926 490813
rect 238050 490873 238084 490889
rect 238050 490797 238084 490813
rect 238168 490873 238202 490889
rect 238168 490797 238202 490813
rect 238326 490873 238360 490889
rect 238326 490797 238360 490813
rect 238444 490873 238478 490889
rect 238444 490797 238478 490813
rect 238602 490873 238636 490889
rect 238602 490797 238636 490813
rect 238720 490873 238754 490889
rect 238720 490797 238754 490813
rect 238878 490873 238912 490889
rect 238878 490797 238912 490813
rect 238996 490873 239030 490889
rect 238996 490797 239030 490813
rect 239154 490873 239188 490889
rect 239154 490797 239188 490813
rect 239272 490873 239306 490889
rect 239272 490797 239306 490813
rect 239430 490873 239464 490889
rect 239430 490797 239464 490813
rect 239548 490873 239582 490889
rect 239548 490797 239582 490813
rect 239706 490873 239740 490889
rect 239706 490797 239740 490813
rect 239824 490873 239858 490889
rect 239824 490797 239858 490813
rect 239982 490873 240016 490889
rect 239982 490797 240016 490813
rect 240100 490873 240134 490889
rect 240100 490797 240134 490813
rect 240258 490873 240292 490889
rect 240258 490797 240292 490813
rect 240376 490873 240410 490889
rect 240376 490797 240410 490813
rect 240534 490873 240568 490889
rect 240534 490797 240568 490813
rect 240652 490873 240686 490889
rect 240652 490797 240686 490813
rect 240810 490873 240844 490889
rect 240810 490797 240844 490813
rect 240928 490873 240962 490889
rect 240928 490797 240962 490813
rect 241086 490873 241120 490889
rect 241086 490797 241120 490813
rect 241204 490873 241238 490889
rect 241204 490797 241238 490813
rect 241362 490873 241396 490889
rect 241362 490797 241396 490813
rect 241480 490873 241514 490889
rect 241480 490797 241514 490813
rect 241638 490873 241672 490889
rect 241638 490797 241672 490813
rect 241756 490873 241790 490889
rect 241756 490797 241790 490813
rect 241914 490873 241948 490889
rect 241914 490797 241948 490813
rect 242032 490873 242066 490889
rect 242032 490797 242066 490813
rect 242190 490873 242224 490889
rect 242190 490797 242224 490813
rect 242308 490873 242342 490889
rect 242308 490797 242342 490813
rect 242466 490873 242500 490889
rect 242466 490797 242500 490813
rect 242584 490873 242618 490889
rect 242584 490797 242618 490813
rect 242742 490873 242776 490889
rect 242742 490797 242776 490813
rect 242860 490873 242894 490889
rect 242860 490797 242894 490813
rect 243018 490873 243052 490889
rect 243018 490797 243052 490813
rect 243136 490873 243170 490889
rect 243136 490797 243170 490813
rect 243294 490873 243328 490889
rect 243294 490797 243328 490813
rect 243412 490873 243446 490889
rect 243412 490797 243446 490813
rect 243570 490873 243604 490889
rect 243570 490797 243604 490813
rect 243688 490873 243722 490889
rect 243688 490797 243722 490813
rect 243846 490873 243880 490889
rect 243846 490797 243880 490813
rect 243964 490873 243998 490889
rect 243964 490797 243998 490813
rect 244122 490873 244156 490889
rect 244122 490797 244156 490813
rect 244240 490873 244274 490889
rect 244240 490797 244274 490813
rect 244398 490873 244432 490889
rect 244398 490797 244432 490813
rect 244516 490873 244550 490889
rect 244516 490797 244550 490813
rect 244674 490873 244708 490889
rect 244674 490797 244708 490813
rect 244792 490873 244826 490889
rect 244792 490797 244826 490813
rect 244950 490873 244984 490889
rect 244950 490797 244984 490813
rect 245068 490873 245102 490889
rect 245068 490797 245102 490813
rect 245226 490873 245260 490889
rect 245226 490797 245260 490813
rect 245344 490873 245378 490889
rect 245344 490797 245378 490813
rect 245502 490873 245536 490889
rect 245502 490797 245536 490813
rect 245620 490873 245654 490889
rect 245620 490797 245654 490813
rect 245778 490873 245812 490889
rect 245778 490797 245812 490813
rect 245896 490873 245930 490889
rect 245896 490797 245930 490813
rect 246054 490873 246088 490889
rect 246054 490797 246088 490813
rect 246172 490873 246206 490889
rect 246172 490797 246206 490813
rect 246330 490873 246364 490889
rect 246330 490797 246364 490813
rect 246448 490873 246482 490889
rect 246448 490797 246482 490813
rect 246606 490873 246640 490889
rect 246606 490797 246640 490813
rect 232694 490729 232710 490763
rect 232778 490760 232794 490763
rect 232778 490729 232802 490760
rect 232970 490729 232986 490763
rect 233054 490729 233070 490763
rect 233246 490759 233262 490763
rect 233243 490729 233262 490759
rect 233330 490729 233346 490763
rect 233522 490755 233538 490763
rect 233519 490729 233538 490755
rect 233606 490729 233622 490763
rect 233798 490749 233814 490763
rect 233797 490729 233814 490749
rect 233882 490729 233898 490763
rect 234074 490745 234090 490763
rect 234073 490729 234090 490745
rect 234158 490729 234174 490763
rect 234350 490747 234366 490763
rect 234347 490729 234366 490747
rect 234434 490729 234450 490763
rect 234626 490745 234642 490763
rect 234625 490729 234642 490745
rect 234710 490729 234726 490763
rect 234902 490729 234918 490763
rect 234986 490729 235002 490763
rect 235178 490745 235194 490763
rect 235177 490729 235194 490745
rect 235262 490729 235278 490763
rect 235454 490729 235470 490763
rect 235538 490729 235554 490763
rect 235730 490755 235746 490763
rect 235727 490739 235746 490755
rect 235726 490729 235746 490739
rect 235814 490729 235830 490763
rect 236006 490755 236022 490763
rect 236003 490729 236022 490755
rect 236090 490729 236106 490763
rect 236282 490729 236298 490763
rect 236366 490729 236382 490763
rect 236558 490749 236574 490763
rect 236551 490729 236574 490749
rect 236642 490729 236658 490763
rect 236834 490729 236850 490763
rect 236918 490729 236934 490763
rect 237110 490749 237126 490763
rect 237109 490729 237126 490749
rect 237194 490729 237210 490763
rect 237386 490745 237402 490763
rect 237385 490729 237402 490745
rect 237470 490729 237486 490763
rect 237662 490753 237678 490763
rect 237659 490729 237678 490753
rect 237746 490729 237762 490763
rect 237938 490745 237954 490763
rect 237937 490729 237954 490745
rect 238022 490729 238038 490763
rect 238214 490747 238230 490763
rect 238207 490729 238230 490747
rect 238298 490729 238314 490763
rect 238490 490753 238506 490763
rect 238483 490729 238506 490753
rect 238574 490729 238590 490763
rect 238766 490759 238782 490763
rect 238765 490729 238782 490759
rect 238850 490729 238866 490763
rect 239042 490755 239058 490763
rect 239041 490729 239058 490755
rect 239126 490729 239142 490763
rect 239318 490755 239334 490763
rect 239315 490729 239334 490755
rect 239402 490729 239418 490763
rect 239594 490755 239610 490763
rect 239587 490729 239610 490755
rect 239678 490729 239694 490763
rect 239870 490755 239886 490763
rect 239869 490729 239886 490755
rect 239954 490729 239970 490763
rect 240146 490729 240162 490763
rect 240230 490729 240246 490763
rect 240422 490749 240438 490763
rect 240421 490729 240438 490749
rect 240506 490729 240522 490763
rect 240698 490729 240714 490763
rect 240782 490729 240798 490763
rect 240974 490729 240990 490763
rect 241058 490729 241074 490763
rect 241250 490741 241266 490763
rect 241243 490729 241266 490741
rect 241334 490729 241350 490763
rect 241526 490737 241542 490763
rect 241525 490729 241542 490737
rect 241610 490729 241626 490763
rect 241802 490729 241818 490763
rect 241886 490729 241902 490763
rect 242078 490737 242094 490763
rect 242077 490729 242094 490737
rect 242162 490729 242178 490763
rect 242354 490737 242370 490763
rect 242353 490729 242370 490737
rect 242438 490729 242454 490763
rect 242630 490753 242646 490763
rect 242623 490729 242646 490753
rect 242714 490729 242730 490763
rect 242906 490745 242922 490763
rect 242901 490729 242922 490745
rect 242990 490729 243006 490763
rect 243182 490729 243198 490763
rect 243266 490729 243282 490763
rect 243458 490729 243474 490763
rect 243542 490745 243558 490763
rect 243734 490749 243750 490763
rect 243542 490729 243563 490745
rect 232700 490520 232802 490729
rect 232971 490520 233069 490729
rect 233243 490520 233341 490729
rect 233519 490520 233617 490729
rect 233797 490520 233895 490729
rect 234073 490520 234171 490729
rect 234347 490520 234445 490729
rect 234625 490520 234723 490729
rect 234903 490520 235001 490729
rect 235177 490520 235275 490729
rect 235455 490520 235553 490729
rect 235726 490520 235826 490729
rect 236003 490520 236101 490729
rect 236283 490520 236381 490729
rect 236551 490520 236649 490729
rect 236835 490520 236933 490729
rect 237109 490520 237207 490729
rect 237385 490520 237483 490729
rect 237659 490520 237757 490729
rect 237937 490520 238035 490729
rect 238207 490520 238305 490729
rect 238483 490520 238581 490729
rect 238765 490520 238863 490729
rect 239041 490520 239139 490729
rect 239315 490714 239413 490729
rect 239587 490520 239685 490729
rect 239869 490520 239967 490729
rect 240147 490520 240245 490729
rect 240421 490520 240519 490729
rect 240699 490520 240797 490729
rect 240975 490520 241073 490729
rect 241243 490520 241341 490729
rect 241525 490520 241623 490729
rect 241803 490520 241901 490729
rect 242077 490520 242175 490729
rect 242353 490520 242451 490729
rect 242623 490520 242721 490729
rect 242901 490520 242999 490729
rect 243183 490520 243281 490729
rect 243465 490520 243563 490729
rect 243733 490729 243750 490749
rect 243818 490729 243834 490763
rect 244010 490749 244026 490763
rect 244009 490729 244026 490749
rect 244094 490729 244110 490763
rect 244286 490749 244302 490763
rect 244279 490729 244302 490749
rect 244370 490729 244386 490763
rect 244562 490755 244578 490763
rect 244557 490729 244578 490755
rect 244646 490729 244662 490763
rect 244838 490729 244854 490763
rect 244922 490729 244938 490763
rect 245114 490729 245130 490763
rect 245198 490755 245214 490763
rect 245198 490729 245217 490755
rect 245390 490753 245406 490763
rect 243733 490520 243831 490729
rect 244009 490520 244107 490729
rect 244279 490520 244377 490729
rect 244557 490520 244655 490729
rect 244839 490520 244937 490729
rect 245119 490520 245217 490729
rect 245385 490729 245406 490753
rect 245474 490729 245490 490763
rect 245666 490747 245682 490763
rect 245661 490729 245682 490747
rect 245750 490729 245766 490763
rect 245942 490753 245958 490763
rect 245941 490729 245958 490753
rect 246026 490729 246042 490763
rect 246218 490729 246234 490763
rect 246302 490753 246318 490763
rect 246302 490729 246323 490753
rect 246494 490729 246510 490763
rect 246578 490757 246594 490763
rect 246578 490729 246601 490757
rect 245385 490520 245483 490729
rect 245661 490520 245759 490729
rect 245941 490520 246039 490729
rect 246225 490520 246323 490729
rect 246503 490520 246601 490729
rect 246740 490671 246774 490687
rect 247092 490520 247190 491144
rect 232697 490489 247190 490520
rect 232697 490433 236703 490489
rect 236781 490433 247190 490489
rect 232697 490422 247190 490433
rect 323888 372598 323968 372608
rect 323888 372556 323904 372598
rect 323958 372556 323968 372598
rect 323888 372231 323968 372556
rect 324161 372488 338373 372515
rect 324160 372417 338373 372488
rect 324160 372231 324258 372417
rect 324436 372231 324534 372417
rect 324710 372231 324808 372417
rect 324988 372231 325086 372417
rect 325260 372231 325358 372417
rect 325538 372231 325636 372417
rect 325816 372231 325914 372417
rect 326094 372231 326192 372417
rect 326368 372231 326466 372417
rect 326644 372231 326742 372417
rect 326920 372231 327018 372417
rect 327198 372231 327296 372417
rect 327474 372231 327572 372417
rect 327746 372231 327844 372417
rect 328024 372231 328122 372417
rect 328296 372231 328394 372417
rect 328574 372231 328672 372417
rect 328850 372231 328948 372417
rect 323877 372197 323893 372231
rect 323961 372197 323977 372231
rect 324153 372197 324169 372231
rect 324237 372206 324258 372231
rect 324237 372197 324253 372206
rect 324429 372197 324445 372231
rect 324513 372208 324534 372231
rect 324513 372197 324529 372208
rect 324705 372197 324721 372231
rect 324789 372204 324808 372231
rect 324789 372197 324805 372204
rect 324981 372197 324997 372231
rect 325065 372204 325086 372231
rect 325065 372197 325081 372204
rect 325257 372197 325273 372231
rect 325341 372206 325358 372231
rect 325341 372197 325357 372206
rect 325533 372197 325549 372231
rect 325617 372204 325636 372231
rect 325617 372197 325633 372204
rect 325809 372197 325825 372231
rect 325893 372204 325914 372231
rect 325893 372197 325909 372204
rect 326085 372197 326101 372231
rect 326169 372208 326192 372231
rect 326169 372197 326185 372208
rect 326361 372197 326377 372231
rect 326445 372204 326466 372231
rect 326445 372197 326461 372204
rect 326637 372197 326653 372231
rect 326721 372208 326742 372231
rect 326721 372197 326737 372208
rect 326913 372197 326929 372231
rect 326997 372208 327018 372231
rect 326997 372197 327013 372208
rect 327189 372197 327205 372231
rect 327273 372210 327296 372231
rect 327273 372197 327289 372210
rect 327465 372197 327481 372231
rect 327549 372200 327572 372231
rect 327549 372197 327565 372200
rect 327741 372197 327757 372231
rect 327825 372204 327844 372231
rect 327825 372197 327841 372204
rect 328017 372197 328033 372231
rect 328101 372204 328122 372231
rect 328101 372197 328117 372204
rect 328293 372197 328309 372231
rect 328377 372197 328394 372231
rect 328569 372197 328585 372231
rect 328653 372204 328672 372231
rect 328653 372197 328669 372204
rect 328845 372197 328861 372231
rect 328929 372204 328948 372231
rect 329120 372231 329218 372417
rect 329406 372231 329504 372417
rect 329678 372231 329776 372417
rect 329958 372231 330056 372417
rect 330232 372231 330330 372417
rect 330508 372231 330606 372417
rect 330784 372231 330882 372417
rect 331060 372231 331158 372417
rect 331336 372231 331434 372417
rect 331612 372231 331710 372417
rect 331888 372231 331986 372417
rect 332164 372231 332262 372417
rect 332442 372231 332540 372417
rect 332718 372231 332816 372417
rect 332990 372231 333088 372417
rect 333268 372231 333366 372417
rect 333544 372231 333642 372417
rect 333822 372231 333920 372417
rect 334096 372231 334194 372417
rect 334372 372231 334470 372417
rect 334650 372231 334748 372417
rect 334926 372231 335024 372417
rect 335202 372231 335300 372417
rect 335478 372231 335576 372417
rect 335754 372231 335852 372417
rect 336028 372231 336126 372417
rect 336308 372231 336406 372417
rect 336584 372231 336682 372417
rect 336856 372231 336954 372417
rect 337132 372231 337230 372417
rect 337402 372231 337500 372417
rect 337694 372231 337792 372417
rect 328929 372197 328945 372204
rect 329120 372202 329137 372231
rect 329121 372197 329137 372202
rect 329205 372197 329221 372231
rect 329397 372197 329413 372231
rect 329481 372200 329504 372231
rect 329481 372197 329497 372200
rect 329673 372197 329689 372231
rect 329757 372200 329776 372231
rect 329757 372197 329773 372200
rect 329949 372197 329965 372231
rect 330033 372200 330056 372231
rect 330033 372197 330049 372200
rect 330225 372197 330241 372231
rect 330309 372200 330330 372231
rect 330309 372197 330325 372200
rect 330501 372197 330517 372231
rect 330585 372202 330606 372231
rect 330585 372197 330601 372202
rect 330777 372197 330793 372231
rect 330861 372200 330882 372231
rect 330861 372197 330877 372200
rect 331053 372197 331069 372231
rect 331137 372202 331158 372231
rect 331137 372197 331153 372202
rect 331329 372197 331345 372231
rect 331413 372202 331434 372231
rect 331413 372197 331429 372202
rect 331605 372197 331621 372231
rect 331689 372204 331710 372231
rect 331689 372197 331705 372204
rect 331881 372197 331897 372231
rect 331965 372202 331986 372231
rect 331965 372197 331981 372202
rect 332157 372197 332173 372231
rect 332241 372202 332262 372231
rect 332241 372197 332257 372202
rect 332433 372197 332449 372231
rect 332517 372202 332540 372231
rect 332517 372197 332533 372202
rect 332709 372197 332725 372231
rect 332793 372202 332816 372231
rect 332793 372197 332809 372202
rect 332985 372197 333001 372231
rect 333069 372200 333088 372231
rect 333069 372197 333085 372200
rect 333261 372197 333277 372231
rect 333345 372200 333366 372231
rect 333345 372197 333361 372200
rect 333537 372197 333553 372231
rect 333621 372204 333642 372231
rect 333621 372197 333637 372204
rect 333813 372197 333829 372231
rect 333897 372206 333920 372231
rect 333897 372197 333913 372206
rect 334089 372197 334105 372231
rect 334173 372202 334194 372231
rect 334173 372197 334189 372202
rect 334365 372197 334381 372231
rect 334449 372206 334470 372231
rect 334449 372197 334465 372206
rect 334641 372197 334657 372231
rect 334725 372206 334748 372231
rect 334725 372197 334741 372206
rect 334917 372197 334933 372231
rect 335001 372208 335024 372231
rect 335001 372197 335017 372208
rect 335193 372197 335209 372231
rect 335277 372204 335300 372231
rect 335277 372197 335293 372204
rect 335469 372197 335485 372231
rect 335553 372206 335576 372231
rect 335553 372197 335569 372206
rect 335745 372197 335761 372231
rect 335829 372206 335852 372231
rect 335829 372197 335845 372206
rect 336021 372197 336037 372231
rect 336105 372208 336126 372231
rect 336105 372197 336121 372208
rect 336297 372197 336313 372231
rect 336381 372208 336406 372231
rect 336381 372197 336397 372208
rect 336573 372197 336589 372231
rect 336657 372208 336682 372231
rect 336657 372197 336673 372208
rect 336849 372197 336865 372231
rect 336933 372208 336954 372231
rect 336933 372197 336949 372208
rect 337125 372197 337141 372231
rect 337209 372198 337230 372231
rect 337209 372197 337225 372198
rect 337401 372197 337417 372231
rect 337485 372197 337501 372231
rect 337677 372197 337693 372231
rect 337761 372198 337792 372231
rect 337923 372273 337957 372289
rect 337761 372197 337777 372198
rect 323888 372192 323968 372197
rect 328296 372196 328394 372197
rect 337402 372196 337500 372197
rect 323831 372147 323865 372163
rect 323831 372071 323865 372087
rect 323989 372147 324023 372163
rect 323989 372071 324023 372087
rect 324107 372147 324141 372163
rect 324107 372071 324141 372087
rect 324265 372147 324299 372163
rect 324265 372071 324299 372087
rect 324383 372147 324417 372163
rect 324383 372071 324417 372087
rect 324541 372147 324575 372163
rect 324541 372071 324575 372087
rect 324659 372147 324693 372163
rect 324659 372071 324693 372087
rect 324817 372147 324851 372163
rect 324817 372071 324851 372087
rect 324935 372147 324969 372163
rect 324935 372071 324969 372087
rect 325093 372147 325127 372163
rect 325093 372071 325127 372087
rect 325211 372147 325245 372163
rect 325211 372071 325245 372087
rect 325369 372147 325403 372163
rect 325369 372071 325403 372087
rect 325487 372147 325521 372163
rect 325487 372071 325521 372087
rect 325645 372147 325679 372163
rect 325645 372071 325679 372087
rect 325763 372147 325797 372163
rect 325763 372071 325797 372087
rect 325921 372147 325955 372163
rect 325921 372071 325955 372087
rect 326039 372147 326073 372163
rect 326039 372071 326073 372087
rect 326197 372147 326231 372163
rect 326197 372071 326231 372087
rect 326315 372147 326349 372163
rect 326315 372071 326349 372087
rect 326473 372147 326507 372163
rect 326473 372071 326507 372087
rect 326591 372147 326625 372163
rect 326591 372071 326625 372087
rect 326749 372147 326783 372163
rect 326749 372071 326783 372087
rect 326867 372147 326901 372163
rect 326867 372071 326901 372087
rect 327025 372147 327059 372163
rect 327025 372071 327059 372087
rect 327143 372147 327177 372163
rect 327143 372071 327177 372087
rect 327301 372147 327335 372163
rect 327301 372071 327335 372087
rect 327419 372147 327453 372163
rect 327419 372071 327453 372087
rect 327577 372147 327611 372163
rect 327577 372071 327611 372087
rect 327695 372147 327729 372163
rect 327695 372071 327729 372087
rect 327853 372147 327887 372163
rect 327853 372071 327887 372087
rect 327971 372147 328005 372163
rect 327971 372071 328005 372087
rect 328129 372147 328163 372163
rect 328129 372071 328163 372087
rect 328247 372147 328281 372163
rect 328247 372071 328281 372087
rect 328405 372147 328439 372163
rect 328405 372071 328439 372087
rect 328523 372147 328557 372163
rect 328523 372071 328557 372087
rect 328681 372147 328715 372163
rect 328681 372071 328715 372087
rect 328799 372147 328833 372163
rect 328799 372071 328833 372087
rect 328957 372147 328991 372163
rect 328957 372071 328991 372087
rect 329075 372147 329109 372163
rect 329075 372071 329109 372087
rect 329233 372147 329267 372163
rect 329233 372071 329267 372087
rect 329351 372147 329385 372163
rect 329351 372071 329385 372087
rect 329509 372147 329543 372163
rect 329509 372071 329543 372087
rect 329627 372147 329661 372163
rect 329627 372071 329661 372087
rect 329785 372147 329819 372163
rect 329785 372071 329819 372087
rect 329903 372147 329937 372163
rect 329903 372071 329937 372087
rect 330061 372147 330095 372163
rect 330061 372071 330095 372087
rect 330179 372147 330213 372163
rect 330179 372071 330213 372087
rect 330337 372147 330371 372163
rect 330337 372071 330371 372087
rect 330455 372147 330489 372163
rect 330455 372071 330489 372087
rect 330613 372147 330647 372163
rect 330613 372071 330647 372087
rect 330731 372147 330765 372163
rect 330731 372071 330765 372087
rect 330889 372147 330923 372163
rect 330889 372071 330923 372087
rect 331007 372147 331041 372163
rect 331007 372071 331041 372087
rect 331165 372147 331199 372163
rect 331165 372071 331199 372087
rect 331283 372147 331317 372163
rect 331283 372071 331317 372087
rect 331441 372147 331475 372163
rect 331441 372071 331475 372087
rect 331559 372147 331593 372163
rect 331559 372071 331593 372087
rect 331717 372147 331751 372163
rect 331717 372071 331751 372087
rect 331835 372147 331869 372163
rect 331835 372071 331869 372087
rect 331993 372147 332027 372163
rect 331993 372071 332027 372087
rect 332111 372147 332145 372163
rect 332111 372071 332145 372087
rect 332269 372147 332303 372163
rect 332269 372071 332303 372087
rect 332387 372147 332421 372163
rect 332387 372071 332421 372087
rect 332545 372147 332579 372163
rect 332545 372071 332579 372087
rect 332663 372147 332697 372163
rect 332663 372071 332697 372087
rect 332821 372147 332855 372163
rect 332821 372071 332855 372087
rect 332939 372147 332973 372163
rect 332939 372071 332973 372087
rect 333097 372147 333131 372163
rect 333097 372071 333131 372087
rect 333215 372147 333249 372163
rect 333215 372071 333249 372087
rect 333373 372147 333407 372163
rect 333373 372071 333407 372087
rect 333491 372147 333525 372163
rect 333491 372071 333525 372087
rect 333649 372147 333683 372163
rect 333649 372071 333683 372087
rect 333767 372147 333801 372163
rect 333767 372071 333801 372087
rect 333925 372147 333959 372163
rect 333925 372071 333959 372087
rect 334043 372147 334077 372163
rect 334043 372071 334077 372087
rect 334201 372147 334235 372163
rect 334201 372071 334235 372087
rect 334319 372147 334353 372163
rect 334319 372071 334353 372087
rect 334477 372147 334511 372163
rect 334477 372071 334511 372087
rect 334595 372147 334629 372163
rect 334595 372071 334629 372087
rect 334753 372147 334787 372163
rect 334753 372071 334787 372087
rect 334871 372147 334905 372163
rect 334871 372071 334905 372087
rect 335029 372147 335063 372163
rect 335029 372071 335063 372087
rect 335147 372147 335181 372163
rect 335147 372071 335181 372087
rect 335305 372147 335339 372163
rect 335305 372071 335339 372087
rect 335423 372147 335457 372163
rect 335423 372071 335457 372087
rect 335581 372147 335615 372163
rect 335581 372071 335615 372087
rect 335699 372147 335733 372163
rect 335699 372071 335733 372087
rect 335857 372147 335891 372163
rect 335857 372071 335891 372087
rect 335975 372147 336009 372163
rect 335975 372071 336009 372087
rect 336133 372147 336167 372163
rect 336133 372071 336167 372087
rect 336251 372147 336285 372163
rect 336251 372071 336285 372087
rect 336409 372147 336443 372163
rect 336409 372071 336443 372087
rect 336527 372147 336561 372163
rect 336527 372071 336561 372087
rect 336685 372147 336719 372163
rect 336685 372071 336719 372087
rect 336803 372147 336837 372163
rect 336803 372071 336837 372087
rect 336961 372147 336995 372163
rect 336961 372071 336995 372087
rect 337079 372147 337113 372163
rect 337079 372071 337113 372087
rect 337237 372147 337271 372163
rect 337237 372071 337271 372087
rect 337355 372147 337389 372163
rect 337355 372071 337389 372087
rect 337513 372147 337547 372163
rect 337513 372071 337547 372087
rect 337631 372147 337665 372163
rect 337631 372071 337665 372087
rect 337789 372147 337823 372163
rect 337789 372071 337823 372087
rect 323888 372037 323968 372040
rect 323877 372003 323893 372037
rect 323961 372003 323977 372037
rect 324153 372003 324169 372037
rect 324237 372003 324253 372037
rect 324429 372032 324445 372037
rect 324426 372003 324445 372032
rect 324513 372003 324529 372037
rect 324705 372028 324721 372037
rect 324702 372003 324721 372028
rect 324789 372003 324805 372037
rect 324981 372022 324997 372037
rect 324980 372003 324997 372022
rect 325065 372003 325081 372037
rect 325257 372018 325273 372037
rect 325256 372003 325273 372018
rect 325341 372003 325357 372037
rect 325533 372020 325549 372037
rect 325530 372003 325549 372020
rect 325617 372003 325633 372037
rect 325809 372018 325825 372037
rect 325808 372003 325825 372018
rect 325893 372003 325909 372037
rect 326085 372003 326101 372037
rect 326169 372003 326185 372037
rect 326361 372018 326377 372037
rect 326360 372003 326377 372018
rect 326445 372003 326461 372037
rect 326637 372003 326653 372037
rect 326721 372003 326737 372037
rect 326913 372028 326929 372037
rect 326910 372003 326929 372028
rect 326997 372003 327013 372037
rect 327189 372028 327205 372037
rect 327186 372003 327205 372028
rect 327273 372003 327289 372037
rect 327465 372003 327481 372037
rect 327549 372003 327565 372037
rect 327741 372022 327757 372037
rect 327734 372003 327757 372022
rect 327825 372003 327841 372037
rect 328017 372003 328033 372037
rect 328101 372003 328117 372037
rect 328293 372022 328309 372037
rect 328292 372003 328309 372022
rect 328377 372003 328393 372037
rect 328569 372018 328585 372037
rect 328568 372003 328585 372018
rect 328653 372003 328669 372037
rect 328845 372026 328861 372037
rect 328842 372003 328861 372026
rect 328929 372003 328945 372037
rect 329121 372018 329137 372037
rect 329120 372003 329137 372018
rect 329205 372003 329221 372037
rect 329397 372020 329413 372037
rect 329390 372003 329413 372020
rect 329481 372003 329497 372037
rect 329673 372026 329689 372037
rect 329666 372003 329689 372026
rect 329757 372003 329773 372037
rect 329949 372032 329965 372037
rect 329948 372003 329965 372032
rect 330033 372003 330049 372037
rect 330225 372028 330241 372037
rect 330224 372003 330241 372028
rect 330309 372003 330325 372037
rect 330501 372028 330517 372037
rect 330498 372003 330517 372028
rect 330585 372003 330601 372037
rect 330777 372028 330793 372037
rect 330770 372003 330793 372028
rect 330861 372003 330877 372037
rect 331053 372028 331069 372037
rect 331052 372003 331069 372028
rect 331137 372003 331153 372037
rect 331329 372003 331345 372037
rect 331413 372003 331429 372037
rect 331605 372022 331621 372037
rect 331604 372003 331621 372022
rect 331689 372003 331705 372037
rect 331881 372003 331897 372037
rect 331965 372003 331981 372037
rect 332157 372003 332173 372037
rect 332241 372003 332257 372037
rect 332433 372014 332449 372037
rect 332426 372003 332449 372014
rect 332517 372003 332533 372037
rect 332709 372010 332725 372037
rect 332708 372003 332725 372010
rect 332793 372003 332809 372037
rect 332985 372003 333001 372037
rect 333069 372003 333085 372037
rect 333261 372010 333277 372037
rect 333260 372003 333277 372010
rect 333345 372003 333361 372037
rect 333537 372010 333553 372037
rect 333536 372003 333553 372010
rect 333621 372003 333637 372037
rect 333813 372026 333829 372037
rect 333806 372003 333829 372026
rect 333897 372003 333913 372037
rect 334089 372018 334105 372037
rect 334084 372003 334105 372018
rect 334173 372003 334189 372037
rect 334365 372003 334381 372037
rect 334449 372003 334465 372037
rect 334641 372003 334657 372037
rect 334725 372018 334741 372037
rect 334917 372022 334933 372037
rect 334725 372003 334746 372018
rect 53336 371780 67833 371838
rect 143336 371780 157833 371838
rect 53335 371740 67833 371780
rect 53335 371553 53422 371740
rect 53620 371553 53718 371740
rect 53896 371553 53994 371740
rect 54170 371553 54268 371740
rect 54448 371553 54546 371740
rect 54720 371553 54818 371740
rect 54998 371553 55096 371740
rect 55276 371553 55374 371740
rect 55554 371553 55652 371740
rect 55828 371553 55926 371740
rect 56104 371553 56202 371740
rect 56389 371553 56484 371740
rect 56658 371553 56756 371740
rect 56934 371553 57032 371740
rect 57206 371553 57304 371740
rect 57484 371553 57582 371740
rect 57756 371553 57854 371740
rect 58034 371553 58132 371740
rect 58310 371553 58408 371740
rect 53335 371530 53353 371553
rect 53337 371519 53353 371530
rect 53421 371519 53437 371553
rect 53613 371519 53629 371553
rect 53697 371529 53718 371553
rect 53697 371519 53713 371529
rect 53889 371519 53905 371553
rect 53973 371531 53994 371553
rect 53973 371519 53989 371531
rect 54165 371519 54181 371553
rect 54249 371527 54268 371553
rect 54249 371519 54265 371527
rect 54441 371519 54457 371553
rect 54525 371527 54546 371553
rect 54525 371519 54541 371527
rect 54717 371519 54733 371553
rect 54801 371529 54818 371553
rect 54801 371519 54817 371529
rect 54993 371519 55009 371553
rect 55077 371527 55096 371553
rect 55077 371519 55093 371527
rect 55269 371519 55285 371553
rect 55353 371527 55374 371553
rect 55353 371519 55369 371527
rect 55545 371519 55561 371553
rect 55629 371531 55652 371553
rect 55629 371519 55645 371531
rect 55821 371519 55837 371553
rect 55905 371527 55926 371553
rect 55905 371519 55921 371527
rect 56097 371519 56113 371553
rect 56181 371531 56202 371553
rect 56181 371519 56197 371531
rect 56373 371519 56389 371553
rect 56457 371530 56484 371553
rect 56457 371519 56473 371530
rect 56649 371519 56665 371553
rect 56733 371533 56756 371553
rect 56733 371519 56749 371533
rect 56925 371519 56941 371553
rect 57009 371523 57032 371553
rect 57009 371519 57025 371523
rect 57201 371519 57217 371553
rect 57285 371527 57304 371553
rect 57285 371519 57301 371527
rect 57477 371519 57493 371553
rect 57561 371527 57582 371553
rect 57561 371519 57577 371527
rect 57753 371519 57769 371553
rect 57837 371519 57854 371553
rect 58029 371519 58045 371553
rect 58113 371527 58132 371553
rect 58113 371519 58129 371527
rect 58305 371519 58321 371553
rect 58389 371527 58408 371553
rect 58580 371553 58678 371740
rect 58866 371553 58964 371740
rect 59138 371553 59236 371740
rect 59418 371553 59516 371740
rect 59692 371553 59790 371740
rect 60244 371553 60342 371740
rect 60520 371553 60618 371740
rect 60796 371553 60894 371740
rect 61072 371553 61170 371740
rect 61348 371553 61446 371740
rect 61624 371553 61722 371740
rect 61902 371553 62000 371740
rect 62178 371553 62276 371740
rect 62450 371553 62548 371740
rect 62728 371553 62826 371740
rect 63004 371553 63102 371740
rect 63282 371553 63380 371740
rect 63556 371553 63654 371740
rect 63832 371553 63930 371740
rect 64110 371553 64208 371740
rect 64386 371553 64484 371740
rect 64662 371553 64760 371740
rect 64938 371553 65036 371740
rect 65214 371553 65312 371740
rect 65488 371553 65586 371740
rect 65768 371553 65866 371740
rect 66044 371553 66142 371740
rect 66316 371553 66414 371740
rect 66592 371553 66690 371740
rect 66862 371553 66960 371740
rect 67154 371553 67252 371740
rect 58389 371519 58405 371527
rect 58580 371525 58597 371553
rect 58581 371519 58597 371525
rect 58665 371519 58681 371553
rect 58857 371519 58873 371553
rect 58941 371523 58964 371553
rect 58941 371519 58957 371523
rect 59133 371519 59149 371553
rect 59217 371523 59236 371553
rect 59217 371519 59233 371523
rect 59409 371519 59425 371553
rect 59493 371523 59516 371553
rect 59493 371519 59509 371523
rect 59685 371519 59701 371553
rect 59769 371523 59790 371553
rect 59769 371519 59785 371523
rect 59961 371519 59977 371553
rect 60045 371519 60061 371553
rect 60237 371519 60253 371553
rect 60321 371523 60342 371553
rect 60321 371519 60337 371523
rect 60513 371519 60529 371553
rect 60597 371525 60618 371553
rect 60597 371519 60613 371525
rect 60789 371519 60805 371553
rect 60873 371525 60894 371553
rect 60873 371519 60889 371525
rect 61065 371519 61081 371553
rect 61149 371527 61170 371553
rect 61149 371519 61165 371527
rect 61341 371519 61357 371553
rect 61425 371525 61446 371553
rect 61425 371519 61441 371525
rect 61617 371519 61633 371553
rect 61701 371525 61722 371553
rect 61701 371519 61717 371525
rect 61893 371519 61909 371553
rect 61977 371525 62000 371553
rect 61977 371519 61993 371525
rect 62169 371519 62185 371553
rect 62253 371525 62276 371553
rect 62253 371519 62269 371525
rect 62445 371519 62461 371553
rect 62529 371523 62548 371553
rect 62529 371519 62545 371523
rect 62721 371519 62737 371553
rect 62805 371523 62826 371553
rect 62805 371519 62821 371523
rect 62997 371519 63013 371553
rect 63081 371527 63102 371553
rect 63081 371519 63097 371527
rect 63273 371519 63289 371553
rect 63357 371529 63380 371553
rect 63357 371519 63373 371529
rect 63549 371519 63565 371553
rect 63633 371525 63654 371553
rect 63633 371519 63649 371525
rect 63825 371519 63841 371553
rect 63909 371529 63930 371553
rect 63909 371519 63925 371529
rect 64101 371519 64117 371553
rect 64185 371529 64208 371553
rect 64185 371519 64201 371529
rect 64377 371519 64393 371553
rect 64461 371531 64484 371553
rect 64461 371519 64477 371531
rect 64653 371519 64669 371553
rect 64737 371527 64760 371553
rect 64737 371519 64753 371527
rect 64929 371519 64945 371553
rect 65013 371529 65036 371553
rect 65013 371519 65029 371529
rect 65205 371519 65221 371553
rect 65289 371529 65312 371553
rect 65289 371519 65305 371529
rect 65481 371519 65497 371553
rect 65565 371531 65586 371553
rect 65565 371519 65581 371531
rect 65757 371519 65773 371553
rect 65841 371531 65866 371553
rect 65841 371519 65857 371531
rect 66033 371519 66049 371553
rect 66117 371531 66142 371553
rect 66117 371519 66133 371531
rect 66309 371519 66325 371553
rect 66393 371531 66414 371553
rect 66393 371519 66409 371531
rect 66585 371519 66601 371553
rect 66669 371521 66690 371553
rect 66669 371519 66685 371521
rect 66861 371519 66877 371553
rect 66945 371519 66961 371553
rect 67137 371519 67153 371553
rect 67221 371521 67252 371553
rect 67383 371595 67417 371611
rect 67221 371519 67237 371521
rect 53291 371469 53325 371485
rect 53291 371393 53325 371409
rect 53449 371469 53483 371485
rect 53449 371393 53483 371409
rect 53567 371469 53601 371485
rect 53567 371393 53601 371409
rect 53725 371469 53759 371485
rect 53725 371393 53759 371409
rect 53843 371469 53877 371485
rect 53843 371393 53877 371409
rect 54001 371469 54035 371485
rect 54001 371393 54035 371409
rect 54119 371469 54153 371485
rect 54119 371393 54153 371409
rect 54277 371469 54311 371485
rect 54277 371393 54311 371409
rect 54395 371469 54429 371485
rect 54395 371393 54429 371409
rect 54553 371469 54587 371485
rect 54553 371393 54587 371409
rect 54671 371469 54705 371485
rect 54671 371393 54705 371409
rect 54829 371469 54863 371485
rect 54829 371393 54863 371409
rect 54947 371469 54981 371485
rect 54947 371393 54981 371409
rect 55105 371469 55139 371485
rect 55105 371393 55139 371409
rect 55223 371469 55257 371485
rect 55223 371393 55257 371409
rect 55381 371469 55415 371485
rect 55381 371393 55415 371409
rect 55499 371469 55533 371485
rect 55499 371393 55533 371409
rect 55657 371469 55691 371485
rect 55657 371393 55691 371409
rect 55775 371469 55809 371485
rect 55775 371393 55809 371409
rect 55933 371469 55967 371485
rect 55933 371393 55967 371409
rect 56051 371469 56085 371485
rect 56051 371393 56085 371409
rect 56209 371469 56243 371485
rect 56209 371393 56243 371409
rect 56327 371469 56361 371485
rect 56327 371393 56361 371409
rect 56485 371469 56519 371485
rect 56485 371393 56519 371409
rect 56603 371469 56637 371485
rect 56603 371393 56637 371409
rect 56761 371469 56795 371485
rect 56761 371393 56795 371409
rect 56879 371469 56913 371485
rect 56879 371393 56913 371409
rect 57037 371469 57071 371485
rect 57037 371393 57071 371409
rect 57155 371469 57189 371485
rect 57155 371393 57189 371409
rect 57313 371469 57347 371485
rect 57313 371393 57347 371409
rect 57431 371469 57465 371485
rect 57431 371393 57465 371409
rect 57589 371469 57623 371485
rect 57589 371393 57623 371409
rect 57707 371469 57741 371485
rect 57707 371393 57741 371409
rect 57865 371469 57899 371485
rect 57865 371393 57899 371409
rect 57983 371469 58017 371485
rect 57983 371393 58017 371409
rect 58141 371469 58175 371485
rect 58141 371393 58175 371409
rect 58259 371469 58293 371485
rect 58259 371393 58293 371409
rect 58417 371469 58451 371485
rect 58417 371393 58451 371409
rect 58535 371469 58569 371485
rect 58535 371393 58569 371409
rect 58693 371469 58727 371485
rect 58693 371393 58727 371409
rect 58811 371469 58845 371485
rect 58811 371393 58845 371409
rect 58969 371469 59003 371485
rect 58969 371393 59003 371409
rect 59087 371469 59121 371485
rect 59087 371393 59121 371409
rect 59245 371469 59279 371485
rect 59245 371393 59279 371409
rect 59363 371469 59397 371485
rect 59363 371393 59397 371409
rect 59521 371469 59555 371485
rect 59521 371393 59555 371409
rect 59639 371469 59673 371485
rect 59639 371393 59673 371409
rect 59797 371469 59831 371485
rect 59797 371393 59831 371409
rect 59915 371469 59949 371485
rect 59915 371393 59949 371409
rect 60073 371469 60107 371485
rect 60073 371393 60107 371409
rect 60191 371469 60225 371485
rect 60191 371393 60225 371409
rect 60349 371469 60383 371485
rect 60349 371393 60383 371409
rect 60467 371469 60501 371485
rect 60467 371393 60501 371409
rect 60625 371469 60659 371485
rect 60625 371393 60659 371409
rect 60743 371469 60777 371485
rect 60743 371393 60777 371409
rect 60901 371469 60935 371485
rect 60901 371393 60935 371409
rect 61019 371469 61053 371485
rect 61019 371393 61053 371409
rect 61177 371469 61211 371485
rect 61177 371393 61211 371409
rect 61295 371469 61329 371485
rect 61295 371393 61329 371409
rect 61453 371469 61487 371485
rect 61453 371393 61487 371409
rect 61571 371469 61605 371485
rect 61571 371393 61605 371409
rect 61729 371469 61763 371485
rect 61729 371393 61763 371409
rect 61847 371469 61881 371485
rect 61847 371393 61881 371409
rect 62005 371469 62039 371485
rect 62005 371393 62039 371409
rect 62123 371469 62157 371485
rect 62123 371393 62157 371409
rect 62281 371469 62315 371485
rect 62281 371393 62315 371409
rect 62399 371469 62433 371485
rect 62399 371393 62433 371409
rect 62557 371469 62591 371485
rect 62557 371393 62591 371409
rect 62675 371469 62709 371485
rect 62675 371393 62709 371409
rect 62833 371469 62867 371485
rect 62833 371393 62867 371409
rect 62951 371469 62985 371485
rect 62951 371393 62985 371409
rect 63109 371469 63143 371485
rect 63109 371393 63143 371409
rect 63227 371469 63261 371485
rect 63227 371393 63261 371409
rect 63385 371469 63419 371485
rect 63385 371393 63419 371409
rect 63503 371469 63537 371485
rect 63503 371393 63537 371409
rect 63661 371469 63695 371485
rect 63661 371393 63695 371409
rect 63779 371469 63813 371485
rect 63779 371393 63813 371409
rect 63937 371469 63971 371485
rect 63937 371393 63971 371409
rect 64055 371469 64089 371485
rect 64055 371393 64089 371409
rect 64213 371469 64247 371485
rect 64213 371393 64247 371409
rect 64331 371469 64365 371485
rect 64331 371393 64365 371409
rect 64489 371469 64523 371485
rect 64489 371393 64523 371409
rect 64607 371469 64641 371485
rect 64607 371393 64641 371409
rect 64765 371469 64799 371485
rect 64765 371393 64799 371409
rect 64883 371469 64917 371485
rect 64883 371393 64917 371409
rect 65041 371469 65075 371485
rect 65041 371393 65075 371409
rect 65159 371469 65193 371485
rect 65159 371393 65193 371409
rect 65317 371469 65351 371485
rect 65317 371393 65351 371409
rect 65435 371469 65469 371485
rect 65435 371393 65469 371409
rect 65593 371469 65627 371485
rect 65593 371393 65627 371409
rect 65711 371469 65745 371485
rect 65711 371393 65745 371409
rect 65869 371469 65903 371485
rect 65869 371393 65903 371409
rect 65987 371469 66021 371485
rect 65987 371393 66021 371409
rect 66145 371469 66179 371485
rect 66145 371393 66179 371409
rect 66263 371469 66297 371485
rect 66263 371393 66297 371409
rect 66421 371469 66455 371485
rect 66421 371393 66455 371409
rect 66539 371469 66573 371485
rect 66539 371393 66573 371409
rect 66697 371469 66731 371485
rect 66697 371393 66731 371409
rect 66815 371469 66849 371485
rect 66815 371393 66849 371409
rect 66973 371469 67007 371485
rect 66973 371393 67007 371409
rect 67091 371469 67125 371485
rect 67091 371393 67125 371409
rect 67249 371469 67283 371485
rect 67249 371393 67283 371409
rect 53337 371325 53353 371359
rect 53421 371356 53437 371359
rect 53421 371325 53445 371356
rect 53613 371325 53629 371359
rect 53697 371325 53713 371359
rect 53889 371355 53905 371359
rect 53886 371325 53905 371355
rect 53973 371325 53989 371359
rect 54165 371351 54181 371359
rect 54162 371325 54181 371351
rect 54249 371325 54265 371359
rect 54441 371345 54457 371359
rect 54440 371325 54457 371345
rect 54525 371325 54541 371359
rect 54717 371341 54733 371359
rect 54716 371325 54733 371341
rect 54801 371325 54817 371359
rect 54993 371343 55009 371359
rect 54990 371325 55009 371343
rect 55077 371325 55093 371359
rect 55269 371341 55285 371359
rect 55268 371325 55285 371341
rect 55353 371325 55369 371359
rect 55545 371325 55561 371359
rect 55629 371325 55645 371359
rect 55821 371341 55837 371359
rect 55820 371325 55837 371341
rect 55905 371325 55921 371359
rect 56097 371325 56113 371359
rect 56181 371325 56197 371359
rect 56373 371351 56389 371359
rect 56370 371335 56389 371351
rect 56369 371325 56389 371335
rect 56457 371325 56473 371359
rect 56649 371351 56665 371359
rect 56646 371325 56665 371351
rect 56733 371325 56749 371359
rect 56925 371325 56941 371359
rect 57009 371325 57025 371359
rect 57201 371345 57217 371359
rect 57194 371325 57217 371345
rect 57285 371325 57301 371359
rect 57477 371325 57493 371359
rect 57561 371325 57577 371359
rect 57753 371345 57769 371359
rect 57752 371325 57769 371345
rect 57837 371325 57853 371359
rect 58029 371341 58045 371359
rect 58028 371325 58045 371341
rect 58113 371325 58129 371359
rect 58305 371349 58321 371359
rect 58302 371325 58321 371349
rect 58389 371325 58405 371359
rect 58581 371341 58597 371359
rect 58580 371325 58597 371341
rect 58665 371325 58681 371359
rect 58857 371343 58873 371359
rect 58850 371325 58873 371343
rect 58941 371325 58957 371359
rect 59133 371349 59149 371359
rect 59126 371325 59149 371349
rect 59217 371325 59233 371359
rect 59409 371355 59425 371359
rect 59408 371325 59425 371355
rect 59493 371325 59509 371359
rect 59685 371351 59701 371359
rect 59684 371325 59701 371351
rect 59769 371325 59785 371359
rect 59961 371351 59977 371359
rect 59958 371325 59977 371351
rect 60045 371325 60061 371359
rect 60237 371351 60253 371359
rect 60230 371325 60253 371351
rect 60321 371325 60337 371359
rect 60513 371351 60529 371359
rect 60512 371325 60529 371351
rect 60597 371325 60613 371359
rect 60789 371325 60805 371359
rect 60873 371325 60889 371359
rect 61065 371345 61081 371359
rect 61064 371325 61081 371345
rect 61149 371325 61165 371359
rect 61341 371325 61357 371359
rect 61425 371325 61441 371359
rect 61617 371325 61633 371359
rect 61701 371325 61717 371359
rect 61893 371337 61909 371359
rect 61886 371325 61909 371337
rect 61977 371325 61993 371359
rect 62169 371333 62185 371359
rect 62168 371325 62185 371333
rect 62253 371325 62269 371359
rect 62445 371325 62461 371359
rect 62529 371325 62545 371359
rect 62721 371333 62737 371359
rect 62720 371325 62737 371333
rect 62805 371325 62821 371359
rect 62997 371333 63013 371359
rect 62996 371325 63013 371333
rect 63081 371325 63097 371359
rect 63273 371349 63289 371359
rect 63266 371325 63289 371349
rect 63357 371325 63373 371359
rect 63549 371341 63565 371359
rect 63544 371325 63565 371341
rect 63633 371325 63649 371359
rect 63825 371325 63841 371359
rect 63909 371325 63925 371359
rect 64101 371325 64117 371359
rect 64185 371341 64201 371359
rect 64377 371345 64393 371359
rect 64185 371325 64206 371341
rect 53343 371116 53445 371325
rect 53614 371116 53712 371325
rect 53886 371116 53984 371325
rect 54162 371116 54260 371325
rect 54440 371116 54538 371325
rect 54716 371116 54814 371325
rect 54990 371116 55088 371325
rect 55268 371116 55366 371325
rect 55546 371116 55644 371325
rect 55820 371116 55918 371325
rect 56098 371116 56196 371325
rect 56369 371116 56469 371325
rect 56646 371116 56744 371325
rect 56926 371116 57024 371325
rect 57194 371116 57292 371325
rect 57478 371116 57576 371325
rect 57752 371116 57850 371325
rect 58028 371116 58126 371325
rect 58302 371116 58400 371325
rect 58580 371116 58678 371325
rect 58850 371116 58948 371325
rect 59126 371116 59224 371325
rect 59408 371116 59506 371325
rect 59684 371116 59782 371325
rect 59958 371310 60056 371325
rect 60230 371116 60328 371325
rect 60512 371116 60610 371325
rect 60790 371116 60888 371325
rect 61064 371116 61162 371325
rect 61342 371116 61440 371325
rect 61618 371116 61716 371325
rect 61886 371116 61984 371325
rect 62168 371116 62266 371325
rect 62446 371116 62544 371325
rect 62720 371116 62818 371325
rect 62996 371116 63094 371325
rect 63266 371116 63364 371325
rect 63544 371116 63642 371325
rect 63826 371116 63924 371325
rect 64108 371116 64206 371325
rect 64376 371325 64393 371345
rect 64461 371325 64477 371359
rect 64653 371345 64669 371359
rect 64652 371325 64669 371345
rect 64737 371325 64753 371359
rect 64929 371345 64945 371359
rect 64922 371325 64945 371345
rect 65013 371325 65029 371359
rect 65205 371351 65221 371359
rect 65200 371325 65221 371351
rect 65289 371325 65305 371359
rect 65481 371325 65497 371359
rect 65565 371325 65581 371359
rect 65757 371325 65773 371359
rect 65841 371351 65857 371359
rect 65841 371325 65860 371351
rect 66033 371349 66049 371359
rect 64376 371116 64474 371325
rect 64652 371116 64750 371325
rect 64922 371116 65020 371325
rect 65200 371116 65298 371325
rect 65482 371116 65580 371325
rect 65762 371116 65860 371325
rect 66028 371325 66049 371349
rect 66117 371325 66133 371359
rect 66309 371343 66325 371359
rect 66304 371325 66325 371343
rect 66393 371325 66409 371359
rect 66585 371349 66601 371359
rect 66584 371325 66601 371349
rect 66669 371325 66685 371359
rect 66861 371325 66877 371359
rect 66945 371349 66961 371359
rect 66945 371325 66966 371349
rect 67137 371325 67153 371359
rect 67221 371353 67237 371359
rect 67221 371325 67244 371353
rect 66028 371116 66126 371325
rect 66304 371116 66402 371325
rect 66584 371116 66682 371325
rect 66868 371116 66966 371325
rect 67146 371116 67244 371325
rect 67383 371267 67417 371283
rect 67735 371116 67833 371740
rect 143335 371740 157833 371780
rect 143335 371553 143422 371740
rect 143620 371553 143718 371740
rect 143896 371553 143994 371740
rect 144170 371553 144268 371740
rect 144448 371553 144546 371740
rect 144720 371553 144818 371740
rect 144998 371553 145096 371740
rect 145276 371553 145374 371740
rect 145554 371553 145652 371740
rect 145828 371553 145926 371740
rect 146104 371553 146202 371740
rect 146389 371553 146484 371740
rect 146658 371553 146756 371740
rect 146934 371553 147032 371740
rect 147206 371553 147304 371740
rect 147484 371553 147582 371740
rect 147756 371553 147854 371740
rect 148034 371553 148132 371740
rect 148310 371553 148408 371740
rect 143335 371530 143353 371553
rect 143337 371519 143353 371530
rect 143421 371519 143437 371553
rect 143613 371519 143629 371553
rect 143697 371529 143718 371553
rect 143697 371519 143713 371529
rect 143889 371519 143905 371553
rect 143973 371531 143994 371553
rect 143973 371519 143989 371531
rect 144165 371519 144181 371553
rect 144249 371527 144268 371553
rect 144249 371519 144265 371527
rect 144441 371519 144457 371553
rect 144525 371527 144546 371553
rect 144525 371519 144541 371527
rect 144717 371519 144733 371553
rect 144801 371529 144818 371553
rect 144801 371519 144817 371529
rect 144993 371519 145009 371553
rect 145077 371527 145096 371553
rect 145077 371519 145093 371527
rect 145269 371519 145285 371553
rect 145353 371527 145374 371553
rect 145353 371519 145369 371527
rect 145545 371519 145561 371553
rect 145629 371531 145652 371553
rect 145629 371519 145645 371531
rect 145821 371519 145837 371553
rect 145905 371527 145926 371553
rect 145905 371519 145921 371527
rect 146097 371519 146113 371553
rect 146181 371531 146202 371553
rect 146181 371519 146197 371531
rect 146373 371519 146389 371553
rect 146457 371530 146484 371553
rect 146457 371519 146473 371530
rect 146649 371519 146665 371553
rect 146733 371533 146756 371553
rect 146733 371519 146749 371533
rect 146925 371519 146941 371553
rect 147009 371523 147032 371553
rect 147009 371519 147025 371523
rect 147201 371519 147217 371553
rect 147285 371527 147304 371553
rect 147285 371519 147301 371527
rect 147477 371519 147493 371553
rect 147561 371527 147582 371553
rect 147561 371519 147577 371527
rect 147753 371519 147769 371553
rect 147837 371519 147854 371553
rect 148029 371519 148045 371553
rect 148113 371527 148132 371553
rect 148113 371519 148129 371527
rect 148305 371519 148321 371553
rect 148389 371527 148408 371553
rect 148580 371553 148678 371740
rect 148866 371553 148964 371740
rect 149138 371553 149236 371740
rect 149418 371553 149516 371740
rect 149692 371553 149790 371740
rect 150244 371553 150342 371740
rect 150520 371553 150618 371740
rect 150796 371553 150894 371740
rect 151072 371553 151170 371740
rect 151348 371553 151446 371740
rect 151624 371553 151722 371740
rect 151902 371553 152000 371740
rect 152178 371553 152276 371740
rect 152450 371553 152548 371740
rect 152728 371553 152826 371740
rect 153004 371553 153102 371740
rect 153282 371553 153380 371740
rect 153556 371553 153654 371740
rect 153832 371553 153930 371740
rect 154110 371553 154208 371740
rect 154386 371553 154484 371740
rect 154662 371553 154760 371740
rect 154938 371553 155036 371740
rect 155214 371553 155312 371740
rect 155488 371553 155586 371740
rect 155768 371553 155866 371740
rect 156044 371553 156142 371740
rect 156316 371553 156414 371740
rect 156592 371553 156690 371740
rect 156862 371553 156960 371740
rect 157154 371553 157252 371740
rect 148389 371519 148405 371527
rect 148580 371525 148597 371553
rect 148581 371519 148597 371525
rect 148665 371519 148681 371553
rect 148857 371519 148873 371553
rect 148941 371523 148964 371553
rect 148941 371519 148957 371523
rect 149133 371519 149149 371553
rect 149217 371523 149236 371553
rect 149217 371519 149233 371523
rect 149409 371519 149425 371553
rect 149493 371523 149516 371553
rect 149493 371519 149509 371523
rect 149685 371519 149701 371553
rect 149769 371523 149790 371553
rect 149769 371519 149785 371523
rect 149961 371519 149977 371553
rect 150045 371519 150061 371553
rect 150237 371519 150253 371553
rect 150321 371523 150342 371553
rect 150321 371519 150337 371523
rect 150513 371519 150529 371553
rect 150597 371525 150618 371553
rect 150597 371519 150613 371525
rect 150789 371519 150805 371553
rect 150873 371525 150894 371553
rect 150873 371519 150889 371525
rect 151065 371519 151081 371553
rect 151149 371527 151170 371553
rect 151149 371519 151165 371527
rect 151341 371519 151357 371553
rect 151425 371525 151446 371553
rect 151425 371519 151441 371525
rect 151617 371519 151633 371553
rect 151701 371525 151722 371553
rect 151701 371519 151717 371525
rect 151893 371519 151909 371553
rect 151977 371525 152000 371553
rect 151977 371519 151993 371525
rect 152169 371519 152185 371553
rect 152253 371525 152276 371553
rect 152253 371519 152269 371525
rect 152445 371519 152461 371553
rect 152529 371523 152548 371553
rect 152529 371519 152545 371523
rect 152721 371519 152737 371553
rect 152805 371523 152826 371553
rect 152805 371519 152821 371523
rect 152997 371519 153013 371553
rect 153081 371527 153102 371553
rect 153081 371519 153097 371527
rect 153273 371519 153289 371553
rect 153357 371529 153380 371553
rect 153357 371519 153373 371529
rect 153549 371519 153565 371553
rect 153633 371525 153654 371553
rect 153633 371519 153649 371525
rect 153825 371519 153841 371553
rect 153909 371529 153930 371553
rect 153909 371519 153925 371529
rect 154101 371519 154117 371553
rect 154185 371529 154208 371553
rect 154185 371519 154201 371529
rect 154377 371519 154393 371553
rect 154461 371531 154484 371553
rect 154461 371519 154477 371531
rect 154653 371519 154669 371553
rect 154737 371527 154760 371553
rect 154737 371519 154753 371527
rect 154929 371519 154945 371553
rect 155013 371529 155036 371553
rect 155013 371519 155029 371529
rect 155205 371519 155221 371553
rect 155289 371529 155312 371553
rect 155289 371519 155305 371529
rect 155481 371519 155497 371553
rect 155565 371531 155586 371553
rect 155565 371519 155581 371531
rect 155757 371519 155773 371553
rect 155841 371531 155866 371553
rect 155841 371519 155857 371531
rect 156033 371519 156049 371553
rect 156117 371531 156142 371553
rect 156117 371519 156133 371531
rect 156309 371519 156325 371553
rect 156393 371531 156414 371553
rect 156393 371519 156409 371531
rect 156585 371519 156601 371553
rect 156669 371521 156690 371553
rect 156669 371519 156685 371521
rect 156861 371519 156877 371553
rect 156945 371519 156961 371553
rect 157137 371519 157153 371553
rect 157221 371521 157252 371553
rect 157383 371595 157417 371611
rect 157221 371519 157237 371521
rect 143291 371469 143325 371485
rect 143291 371393 143325 371409
rect 143449 371469 143483 371485
rect 143449 371393 143483 371409
rect 143567 371469 143601 371485
rect 143567 371393 143601 371409
rect 143725 371469 143759 371485
rect 143725 371393 143759 371409
rect 143843 371469 143877 371485
rect 143843 371393 143877 371409
rect 144001 371469 144035 371485
rect 144001 371393 144035 371409
rect 144119 371469 144153 371485
rect 144119 371393 144153 371409
rect 144277 371469 144311 371485
rect 144277 371393 144311 371409
rect 144395 371469 144429 371485
rect 144395 371393 144429 371409
rect 144553 371469 144587 371485
rect 144553 371393 144587 371409
rect 144671 371469 144705 371485
rect 144671 371393 144705 371409
rect 144829 371469 144863 371485
rect 144829 371393 144863 371409
rect 144947 371469 144981 371485
rect 144947 371393 144981 371409
rect 145105 371469 145139 371485
rect 145105 371393 145139 371409
rect 145223 371469 145257 371485
rect 145223 371393 145257 371409
rect 145381 371469 145415 371485
rect 145381 371393 145415 371409
rect 145499 371469 145533 371485
rect 145499 371393 145533 371409
rect 145657 371469 145691 371485
rect 145657 371393 145691 371409
rect 145775 371469 145809 371485
rect 145775 371393 145809 371409
rect 145933 371469 145967 371485
rect 145933 371393 145967 371409
rect 146051 371469 146085 371485
rect 146051 371393 146085 371409
rect 146209 371469 146243 371485
rect 146209 371393 146243 371409
rect 146327 371469 146361 371485
rect 146327 371393 146361 371409
rect 146485 371469 146519 371485
rect 146485 371393 146519 371409
rect 146603 371469 146637 371485
rect 146603 371393 146637 371409
rect 146761 371469 146795 371485
rect 146761 371393 146795 371409
rect 146879 371469 146913 371485
rect 146879 371393 146913 371409
rect 147037 371469 147071 371485
rect 147037 371393 147071 371409
rect 147155 371469 147189 371485
rect 147155 371393 147189 371409
rect 147313 371469 147347 371485
rect 147313 371393 147347 371409
rect 147431 371469 147465 371485
rect 147431 371393 147465 371409
rect 147589 371469 147623 371485
rect 147589 371393 147623 371409
rect 147707 371469 147741 371485
rect 147707 371393 147741 371409
rect 147865 371469 147899 371485
rect 147865 371393 147899 371409
rect 147983 371469 148017 371485
rect 147983 371393 148017 371409
rect 148141 371469 148175 371485
rect 148141 371393 148175 371409
rect 148259 371469 148293 371485
rect 148259 371393 148293 371409
rect 148417 371469 148451 371485
rect 148417 371393 148451 371409
rect 148535 371469 148569 371485
rect 148535 371393 148569 371409
rect 148693 371469 148727 371485
rect 148693 371393 148727 371409
rect 148811 371469 148845 371485
rect 148811 371393 148845 371409
rect 148969 371469 149003 371485
rect 148969 371393 149003 371409
rect 149087 371469 149121 371485
rect 149087 371393 149121 371409
rect 149245 371469 149279 371485
rect 149245 371393 149279 371409
rect 149363 371469 149397 371485
rect 149363 371393 149397 371409
rect 149521 371469 149555 371485
rect 149521 371393 149555 371409
rect 149639 371469 149673 371485
rect 149639 371393 149673 371409
rect 149797 371469 149831 371485
rect 149797 371393 149831 371409
rect 149915 371469 149949 371485
rect 149915 371393 149949 371409
rect 150073 371469 150107 371485
rect 150073 371393 150107 371409
rect 150191 371469 150225 371485
rect 150191 371393 150225 371409
rect 150349 371469 150383 371485
rect 150349 371393 150383 371409
rect 150467 371469 150501 371485
rect 150467 371393 150501 371409
rect 150625 371469 150659 371485
rect 150625 371393 150659 371409
rect 150743 371469 150777 371485
rect 150743 371393 150777 371409
rect 150901 371469 150935 371485
rect 150901 371393 150935 371409
rect 151019 371469 151053 371485
rect 151019 371393 151053 371409
rect 151177 371469 151211 371485
rect 151177 371393 151211 371409
rect 151295 371469 151329 371485
rect 151295 371393 151329 371409
rect 151453 371469 151487 371485
rect 151453 371393 151487 371409
rect 151571 371469 151605 371485
rect 151571 371393 151605 371409
rect 151729 371469 151763 371485
rect 151729 371393 151763 371409
rect 151847 371469 151881 371485
rect 151847 371393 151881 371409
rect 152005 371469 152039 371485
rect 152005 371393 152039 371409
rect 152123 371469 152157 371485
rect 152123 371393 152157 371409
rect 152281 371469 152315 371485
rect 152281 371393 152315 371409
rect 152399 371469 152433 371485
rect 152399 371393 152433 371409
rect 152557 371469 152591 371485
rect 152557 371393 152591 371409
rect 152675 371469 152709 371485
rect 152675 371393 152709 371409
rect 152833 371469 152867 371485
rect 152833 371393 152867 371409
rect 152951 371469 152985 371485
rect 152951 371393 152985 371409
rect 153109 371469 153143 371485
rect 153109 371393 153143 371409
rect 153227 371469 153261 371485
rect 153227 371393 153261 371409
rect 153385 371469 153419 371485
rect 153385 371393 153419 371409
rect 153503 371469 153537 371485
rect 153503 371393 153537 371409
rect 153661 371469 153695 371485
rect 153661 371393 153695 371409
rect 153779 371469 153813 371485
rect 153779 371393 153813 371409
rect 153937 371469 153971 371485
rect 153937 371393 153971 371409
rect 154055 371469 154089 371485
rect 154055 371393 154089 371409
rect 154213 371469 154247 371485
rect 154213 371393 154247 371409
rect 154331 371469 154365 371485
rect 154331 371393 154365 371409
rect 154489 371469 154523 371485
rect 154489 371393 154523 371409
rect 154607 371469 154641 371485
rect 154607 371393 154641 371409
rect 154765 371469 154799 371485
rect 154765 371393 154799 371409
rect 154883 371469 154917 371485
rect 154883 371393 154917 371409
rect 155041 371469 155075 371485
rect 155041 371393 155075 371409
rect 155159 371469 155193 371485
rect 155159 371393 155193 371409
rect 155317 371469 155351 371485
rect 155317 371393 155351 371409
rect 155435 371469 155469 371485
rect 155435 371393 155469 371409
rect 155593 371469 155627 371485
rect 155593 371393 155627 371409
rect 155711 371469 155745 371485
rect 155711 371393 155745 371409
rect 155869 371469 155903 371485
rect 155869 371393 155903 371409
rect 155987 371469 156021 371485
rect 155987 371393 156021 371409
rect 156145 371469 156179 371485
rect 156145 371393 156179 371409
rect 156263 371469 156297 371485
rect 156263 371393 156297 371409
rect 156421 371469 156455 371485
rect 156421 371393 156455 371409
rect 156539 371469 156573 371485
rect 156539 371393 156573 371409
rect 156697 371469 156731 371485
rect 156697 371393 156731 371409
rect 156815 371469 156849 371485
rect 156815 371393 156849 371409
rect 156973 371469 157007 371485
rect 156973 371393 157007 371409
rect 157091 371469 157125 371485
rect 157091 371393 157125 371409
rect 157249 371469 157283 371485
rect 157249 371393 157283 371409
rect 143337 371325 143353 371359
rect 143421 371356 143437 371359
rect 143421 371325 143445 371356
rect 143613 371325 143629 371359
rect 143697 371325 143713 371359
rect 143889 371355 143905 371359
rect 143886 371325 143905 371355
rect 143973 371325 143989 371359
rect 144165 371351 144181 371359
rect 144162 371325 144181 371351
rect 144249 371325 144265 371359
rect 144441 371345 144457 371359
rect 144440 371325 144457 371345
rect 144525 371325 144541 371359
rect 144717 371341 144733 371359
rect 144716 371325 144733 371341
rect 144801 371325 144817 371359
rect 144993 371343 145009 371359
rect 144990 371325 145009 371343
rect 145077 371325 145093 371359
rect 145269 371341 145285 371359
rect 145268 371325 145285 371341
rect 145353 371325 145369 371359
rect 145545 371325 145561 371359
rect 145629 371325 145645 371359
rect 145821 371341 145837 371359
rect 145820 371325 145837 371341
rect 145905 371325 145921 371359
rect 146097 371325 146113 371359
rect 146181 371325 146197 371359
rect 146373 371351 146389 371359
rect 146370 371335 146389 371351
rect 146369 371325 146389 371335
rect 146457 371325 146473 371359
rect 146649 371351 146665 371359
rect 146646 371325 146665 371351
rect 146733 371325 146749 371359
rect 146925 371325 146941 371359
rect 147009 371325 147025 371359
rect 147201 371345 147217 371359
rect 147194 371325 147217 371345
rect 147285 371325 147301 371359
rect 147477 371325 147493 371359
rect 147561 371325 147577 371359
rect 147753 371345 147769 371359
rect 147752 371325 147769 371345
rect 147837 371325 147853 371359
rect 148029 371341 148045 371359
rect 148028 371325 148045 371341
rect 148113 371325 148129 371359
rect 148305 371349 148321 371359
rect 148302 371325 148321 371349
rect 148389 371325 148405 371359
rect 148581 371341 148597 371359
rect 148580 371325 148597 371341
rect 148665 371325 148681 371359
rect 148857 371343 148873 371359
rect 148850 371325 148873 371343
rect 148941 371325 148957 371359
rect 149133 371349 149149 371359
rect 149126 371325 149149 371349
rect 149217 371325 149233 371359
rect 149409 371355 149425 371359
rect 149408 371325 149425 371355
rect 149493 371325 149509 371359
rect 149685 371351 149701 371359
rect 149684 371325 149701 371351
rect 149769 371325 149785 371359
rect 149961 371351 149977 371359
rect 149958 371325 149977 371351
rect 150045 371325 150061 371359
rect 150237 371351 150253 371359
rect 150230 371325 150253 371351
rect 150321 371325 150337 371359
rect 150513 371351 150529 371359
rect 150512 371325 150529 371351
rect 150597 371325 150613 371359
rect 150789 371325 150805 371359
rect 150873 371325 150889 371359
rect 151065 371345 151081 371359
rect 151064 371325 151081 371345
rect 151149 371325 151165 371359
rect 151341 371325 151357 371359
rect 151425 371325 151441 371359
rect 151617 371325 151633 371359
rect 151701 371325 151717 371359
rect 151893 371337 151909 371359
rect 151886 371325 151909 371337
rect 151977 371325 151993 371359
rect 152169 371333 152185 371359
rect 152168 371325 152185 371333
rect 152253 371325 152269 371359
rect 152445 371325 152461 371359
rect 152529 371325 152545 371359
rect 152721 371333 152737 371359
rect 152720 371325 152737 371333
rect 152805 371325 152821 371359
rect 152997 371333 153013 371359
rect 152996 371325 153013 371333
rect 153081 371325 153097 371359
rect 153273 371349 153289 371359
rect 153266 371325 153289 371349
rect 153357 371325 153373 371359
rect 153549 371341 153565 371359
rect 153544 371325 153565 371341
rect 153633 371325 153649 371359
rect 153825 371325 153841 371359
rect 153909 371325 153925 371359
rect 154101 371325 154117 371359
rect 154185 371341 154201 371359
rect 154377 371345 154393 371359
rect 154185 371325 154206 371341
rect 143343 371116 143445 371325
rect 143614 371116 143712 371325
rect 143886 371116 143984 371325
rect 144162 371116 144260 371325
rect 144440 371116 144538 371325
rect 144716 371116 144814 371325
rect 144990 371116 145088 371325
rect 145268 371116 145366 371325
rect 145546 371116 145644 371325
rect 145820 371116 145918 371325
rect 146098 371116 146196 371325
rect 146369 371116 146469 371325
rect 146646 371116 146744 371325
rect 146926 371116 147024 371325
rect 147194 371116 147292 371325
rect 147478 371116 147576 371325
rect 147752 371116 147850 371325
rect 148028 371116 148126 371325
rect 148302 371116 148400 371325
rect 148580 371116 148678 371325
rect 148850 371116 148948 371325
rect 149126 371116 149224 371325
rect 149408 371116 149506 371325
rect 149684 371116 149782 371325
rect 149958 371310 150056 371325
rect 150230 371116 150328 371325
rect 150512 371116 150610 371325
rect 150790 371116 150888 371325
rect 151064 371116 151162 371325
rect 151342 371116 151440 371325
rect 151618 371116 151716 371325
rect 151886 371116 151984 371325
rect 152168 371116 152266 371325
rect 152446 371116 152544 371325
rect 152720 371116 152818 371325
rect 152996 371116 153094 371325
rect 153266 371116 153364 371325
rect 153544 371116 153642 371325
rect 153826 371116 153924 371325
rect 154108 371116 154206 371325
rect 154376 371325 154393 371345
rect 154461 371325 154477 371359
rect 154653 371345 154669 371359
rect 154652 371325 154669 371345
rect 154737 371325 154753 371359
rect 154929 371345 154945 371359
rect 154922 371325 154945 371345
rect 155013 371325 155029 371359
rect 155205 371351 155221 371359
rect 155200 371325 155221 371351
rect 155289 371325 155305 371359
rect 155481 371325 155497 371359
rect 155565 371325 155581 371359
rect 155757 371325 155773 371359
rect 155841 371351 155857 371359
rect 155841 371325 155860 371351
rect 156033 371349 156049 371359
rect 154376 371116 154474 371325
rect 154652 371116 154750 371325
rect 154922 371116 155020 371325
rect 155200 371116 155298 371325
rect 155482 371116 155580 371325
rect 155762 371116 155860 371325
rect 156028 371325 156049 371349
rect 156117 371325 156133 371359
rect 156309 371343 156325 371359
rect 156304 371325 156325 371343
rect 156393 371325 156409 371359
rect 156585 371349 156601 371359
rect 156584 371325 156601 371349
rect 156669 371325 156685 371359
rect 156861 371325 156877 371359
rect 156945 371349 156961 371359
rect 156945 371325 156966 371349
rect 157137 371325 157153 371359
rect 157221 371353 157237 371359
rect 157221 371325 157244 371353
rect 156028 371116 156126 371325
rect 156304 371116 156402 371325
rect 156584 371116 156682 371325
rect 156868 371116 156966 371325
rect 157146 371116 157244 371325
rect 157383 371267 157417 371283
rect 157735 371116 157833 371740
rect 323888 371686 323968 372003
rect 324154 371793 324252 372003
rect 324426 371793 324524 372003
rect 324702 371793 324800 372003
rect 324980 371793 325078 372003
rect 325256 371793 325354 372003
rect 325530 371793 325628 372003
rect 325808 371793 325906 372003
rect 326086 371793 326184 372003
rect 326360 371793 326458 372003
rect 326638 371793 326736 372003
rect 326910 371793 327008 372003
rect 327186 371793 327284 372003
rect 327466 371793 327564 372003
rect 327734 371793 327832 372003
rect 328018 371793 328116 372003
rect 328292 371793 328390 372003
rect 328568 371793 328666 372003
rect 328842 371793 328940 372003
rect 329120 371793 329218 372003
rect 329390 371793 329488 372003
rect 329666 371793 329764 372003
rect 329948 371793 330046 372003
rect 330224 371793 330322 372003
rect 330498 371793 330596 372003
rect 330770 371793 330868 372003
rect 331052 371793 331150 372003
rect 331330 371793 331428 372003
rect 331604 371793 331702 372003
rect 331882 371793 331980 372003
rect 332158 371793 332256 372003
rect 332426 371793 332524 372003
rect 332708 371793 332806 372003
rect 332986 371793 333084 372003
rect 333260 371793 333358 372003
rect 333536 371793 333634 372003
rect 333806 371793 333904 372003
rect 334084 371793 334182 372003
rect 334366 371793 334464 372003
rect 334648 371793 334746 372003
rect 334916 372003 334933 372022
rect 335001 372003 335017 372037
rect 335193 372022 335209 372037
rect 335192 372003 335209 372022
rect 335277 372003 335293 372037
rect 335469 372022 335485 372037
rect 335462 372003 335485 372022
rect 335553 372003 335569 372037
rect 335745 372028 335761 372037
rect 335740 372003 335761 372028
rect 335829 372003 335845 372037
rect 336021 372003 336037 372037
rect 336105 372003 336121 372037
rect 336297 372003 336313 372037
rect 336381 372028 336397 372037
rect 336381 372003 336400 372028
rect 336573 372026 336589 372037
rect 334916 371793 335014 372003
rect 335192 371793 335290 372003
rect 335462 371793 335560 372003
rect 335740 371793 335838 372003
rect 336022 371793 336120 372003
rect 336302 371793 336400 372003
rect 336568 372003 336589 372026
rect 336657 372003 336673 372037
rect 336849 372020 336865 372037
rect 336844 372003 336865 372020
rect 336933 372003 336949 372037
rect 337125 372026 337141 372037
rect 337124 372003 337141 372026
rect 337209 372003 337225 372037
rect 337401 372003 337417 372037
rect 337485 372026 337501 372037
rect 337485 372003 337506 372026
rect 337677 372003 337693 372037
rect 337761 372030 337777 372037
rect 337761 372003 337784 372030
rect 336568 371793 336666 372003
rect 336844 371793 336942 372003
rect 337124 371793 337222 372003
rect 337408 371793 337506 372003
rect 337686 371793 337784 372003
rect 337923 371945 337957 371961
rect 338275 371793 338373 372417
rect 324154 371762 338373 371793
rect 324154 371706 327886 371762
rect 327964 371706 338373 371762
rect 324154 371695 338373 371706
rect 418580 371988 421459 371999
rect 418580 371957 421460 371988
rect 323888 371644 323904 371686
rect 323958 371644 323968 371686
rect 323888 371624 323968 371644
rect 418580 371514 418622 371957
rect 418900 371952 421460 371957
rect 418900 371843 418978 371952
rect 419176 371843 419254 371952
rect 419454 371843 419532 371952
rect 419726 371843 419804 371952
rect 420008 371843 420086 371850
rect 420280 371843 420358 371952
rect 420556 371843 420634 371952
rect 420830 371843 420908 371952
rect 421108 371843 421186 371952
rect 421382 371843 421460 371952
rect 421617 371885 421651 371901
rect 418887 371809 418903 371843
rect 418971 371809 418987 371843
rect 419163 371809 419179 371843
rect 419247 371809 419263 371843
rect 419439 371809 419455 371843
rect 419523 371809 419539 371843
rect 419715 371809 419731 371843
rect 419799 371809 419815 371843
rect 419991 371809 420007 371843
rect 420075 371809 420091 371843
rect 420267 371809 420283 371843
rect 420351 371809 420367 371843
rect 420543 371809 420559 371843
rect 420627 371809 420643 371843
rect 420819 371809 420835 371843
rect 420903 371809 420919 371843
rect 421095 371809 421111 371843
rect 421179 371809 421195 371843
rect 421371 371809 421387 371843
rect 421455 371809 421471 371843
rect 418900 371808 418978 371809
rect 419176 371806 419254 371809
rect 419454 371808 419532 371809
rect 419726 371808 419804 371809
rect 420008 371808 420086 371809
rect 420280 371808 420358 371809
rect 420556 371806 420634 371809
rect 420830 371806 420908 371809
rect 421108 371808 421186 371809
rect 421382 371806 421460 371809
rect 418841 371759 418875 371775
rect 418841 371683 418875 371699
rect 418999 371759 419033 371775
rect 418999 371683 419033 371699
rect 419117 371759 419151 371775
rect 419117 371683 419151 371699
rect 419275 371759 419309 371775
rect 419275 371683 419309 371699
rect 419393 371759 419427 371775
rect 419393 371683 419427 371699
rect 419551 371759 419585 371775
rect 419551 371683 419585 371699
rect 419669 371759 419703 371775
rect 419669 371683 419703 371699
rect 419827 371759 419861 371775
rect 419827 371683 419861 371699
rect 419945 371759 419979 371775
rect 419945 371683 419979 371699
rect 420103 371759 420137 371775
rect 420103 371683 420137 371699
rect 420221 371759 420255 371775
rect 420221 371683 420255 371699
rect 420379 371759 420413 371775
rect 420379 371683 420413 371699
rect 420497 371759 420531 371775
rect 420497 371683 420531 371699
rect 420655 371759 420689 371775
rect 420655 371683 420689 371699
rect 420773 371759 420807 371775
rect 420773 371683 420807 371699
rect 420931 371759 420965 371775
rect 420931 371683 420965 371699
rect 421049 371759 421083 371775
rect 421049 371683 421083 371699
rect 421207 371759 421241 371775
rect 421207 371683 421241 371699
rect 421325 371759 421359 371775
rect 421325 371683 421359 371699
rect 421483 371759 421517 371775
rect 421483 371683 421517 371699
rect 418904 371649 418982 371650
rect 419730 371649 419808 371650
rect 420006 371649 420084 371650
rect 420278 371649 420356 371652
rect 420556 371649 420634 371650
rect 420834 371649 420912 371652
rect 421110 371649 421188 371652
rect 421386 371649 421464 371654
rect 418887 371615 418903 371649
rect 418971 371615 418987 371649
rect 419163 371615 419179 371649
rect 419247 371615 419263 371649
rect 419439 371615 419455 371649
rect 419523 371615 419539 371649
rect 419715 371615 419731 371649
rect 419799 371615 419815 371649
rect 419991 371615 420007 371649
rect 420075 371615 420091 371649
rect 420267 371615 420283 371649
rect 420351 371615 420367 371649
rect 420543 371615 420559 371649
rect 420627 371615 420643 371649
rect 420819 371615 420835 371649
rect 420903 371615 420919 371649
rect 421095 371615 421111 371649
rect 421179 371615 421195 371649
rect 421371 371615 421387 371649
rect 421455 371615 421471 371649
rect 418904 371514 418982 371615
rect 419178 371514 419256 371615
rect 419454 371514 419532 371615
rect 419730 371514 419808 371615
rect 420006 371608 420084 371615
rect 420278 371514 420356 371615
rect 420556 371514 420634 371615
rect 420834 371514 420912 371615
rect 421110 371514 421188 371615
rect 421386 371514 421464 371615
rect 421617 371557 421651 371573
rect 508707 371582 510075 371618
rect 418580 371472 421466 371514
rect 419544 371334 419660 371472
rect 419544 371290 419566 371334
rect 419638 371290 419660 371334
rect 419544 371264 419660 371290
rect 419602 371258 419660 371264
rect 508707 371246 508743 371582
rect 508907 371515 508977 371582
rect 509175 371515 509245 371582
rect 509723 371515 509793 371582
rect 510005 371515 510075 371582
rect 510236 371557 510270 371573
rect 508886 371481 508902 371515
rect 508970 371481 508986 371515
rect 509162 371481 509178 371515
rect 509246 371481 509262 371515
rect 509438 371481 509454 371515
rect 509522 371481 509538 371515
rect 509714 371481 509730 371515
rect 509798 371481 509814 371515
rect 509990 371481 510006 371515
rect 510074 371481 510090 371515
rect 508907 371476 508977 371481
rect 509175 371476 509245 371481
rect 509723 371474 509793 371481
rect 510005 371476 510075 371481
rect 508840 371431 508874 371447
rect 508840 371355 508874 371371
rect 508998 371431 509032 371447
rect 508998 371355 509032 371371
rect 509116 371431 509150 371447
rect 509116 371355 509150 371371
rect 509274 371431 509308 371447
rect 509274 371355 509308 371371
rect 509392 371431 509426 371447
rect 509392 371355 509426 371371
rect 509550 371431 509584 371447
rect 509550 371355 509584 371371
rect 509668 371431 509702 371447
rect 509668 371355 509702 371371
rect 509826 371431 509860 371447
rect 509826 371355 509860 371371
rect 509944 371431 509978 371447
rect 509944 371355 509978 371371
rect 510102 371431 510136 371447
rect 510102 371355 510136 371371
rect 509721 371321 509817 371322
rect 508886 371287 508902 371321
rect 508970 371287 508986 371321
rect 509162 371287 509178 371321
rect 509246 371287 509262 371321
rect 509438 371287 509454 371321
rect 509522 371287 509538 371321
rect 509714 371287 509730 371321
rect 509798 371287 509817 371321
rect 509990 371287 510006 371321
rect 510074 371287 510090 371321
rect 509165 371246 509259 371287
rect 509721 371250 509817 371287
rect 510011 371260 510075 371287
rect 510011 371250 510073 371260
rect 509719 371246 510073 371250
rect 508707 371244 510073 371246
rect 232693 371184 247190 371242
rect 508707 371210 508923 371244
rect 508961 371210 510073 371244
rect 510236 371229 510270 371245
rect 509719 371208 510073 371210
rect 53340 371085 67833 371116
rect 53340 371029 57346 371085
rect 57424 371029 67833 371085
rect 53340 371018 67833 371029
rect 143340 371085 157833 371116
rect 143340 371029 147346 371085
rect 147424 371029 157833 371085
rect 143340 371018 157833 371029
rect 232692 371144 247190 371184
rect 232692 370957 232779 371144
rect 232977 370957 233075 371144
rect 233253 370957 233351 371144
rect 233527 370957 233625 371144
rect 233805 370957 233903 371144
rect 234077 370957 234175 371144
rect 234355 370957 234453 371144
rect 234633 370957 234731 371144
rect 234911 370957 235009 371144
rect 235185 370957 235283 371144
rect 235461 370957 235559 371144
rect 235746 370957 235841 371144
rect 236015 370957 236113 371144
rect 236291 370957 236389 371144
rect 236563 370957 236661 371144
rect 236841 370957 236939 371144
rect 237113 370957 237211 371144
rect 237391 370957 237489 371144
rect 237667 370957 237765 371144
rect 232692 370934 232710 370957
rect 232694 370923 232710 370934
rect 232778 370923 232794 370957
rect 232970 370923 232986 370957
rect 233054 370933 233075 370957
rect 233054 370923 233070 370933
rect 233246 370923 233262 370957
rect 233330 370935 233351 370957
rect 233330 370923 233346 370935
rect 233522 370923 233538 370957
rect 233606 370931 233625 370957
rect 233606 370923 233622 370931
rect 233798 370923 233814 370957
rect 233882 370931 233903 370957
rect 233882 370923 233898 370931
rect 234074 370923 234090 370957
rect 234158 370933 234175 370957
rect 234158 370923 234174 370933
rect 234350 370923 234366 370957
rect 234434 370931 234453 370957
rect 234434 370923 234450 370931
rect 234626 370923 234642 370957
rect 234710 370931 234731 370957
rect 234710 370923 234726 370931
rect 234902 370923 234918 370957
rect 234986 370935 235009 370957
rect 234986 370923 235002 370935
rect 235178 370923 235194 370957
rect 235262 370931 235283 370957
rect 235262 370923 235278 370931
rect 235454 370923 235470 370957
rect 235538 370935 235559 370957
rect 235538 370923 235554 370935
rect 235730 370923 235746 370957
rect 235814 370934 235841 370957
rect 235814 370923 235830 370934
rect 236006 370923 236022 370957
rect 236090 370937 236113 370957
rect 236090 370923 236106 370937
rect 236282 370923 236298 370957
rect 236366 370927 236389 370957
rect 236366 370923 236382 370927
rect 236558 370923 236574 370957
rect 236642 370931 236661 370957
rect 236642 370923 236658 370931
rect 236834 370923 236850 370957
rect 236918 370931 236939 370957
rect 236918 370923 236934 370931
rect 237110 370923 237126 370957
rect 237194 370923 237211 370957
rect 237386 370923 237402 370957
rect 237470 370931 237489 370957
rect 237470 370923 237486 370931
rect 237662 370923 237678 370957
rect 237746 370931 237765 370957
rect 237937 370957 238035 371144
rect 238223 370957 238321 371144
rect 238495 370957 238593 371144
rect 238775 370957 238873 371144
rect 239049 370957 239147 371144
rect 239601 370957 239699 371144
rect 239877 370957 239975 371144
rect 240153 370957 240251 371144
rect 240429 370957 240527 371144
rect 240705 370957 240803 371144
rect 240981 370957 241079 371144
rect 241259 370957 241357 371144
rect 241535 370957 241633 371144
rect 241807 370957 241905 371144
rect 242085 370957 242183 371144
rect 242361 370957 242459 371144
rect 242639 370957 242737 371144
rect 242913 370957 243011 371144
rect 243189 370957 243287 371144
rect 243467 370957 243565 371144
rect 243743 370957 243841 371144
rect 244019 370957 244117 371144
rect 244295 370957 244393 371144
rect 244571 370957 244669 371144
rect 244845 370957 244943 371144
rect 245125 370957 245223 371144
rect 245401 370957 245499 371144
rect 245673 370957 245771 371144
rect 245949 370957 246047 371144
rect 246219 370957 246317 371144
rect 246511 370957 246609 371144
rect 237746 370923 237762 370931
rect 237937 370929 237954 370957
rect 237938 370923 237954 370929
rect 238022 370923 238038 370957
rect 238214 370923 238230 370957
rect 238298 370927 238321 370957
rect 238298 370923 238314 370927
rect 238490 370923 238506 370957
rect 238574 370927 238593 370957
rect 238574 370923 238590 370927
rect 238766 370923 238782 370957
rect 238850 370927 238873 370957
rect 238850 370923 238866 370927
rect 239042 370923 239058 370957
rect 239126 370927 239147 370957
rect 239126 370923 239142 370927
rect 239318 370923 239334 370957
rect 239402 370923 239418 370957
rect 239594 370923 239610 370957
rect 239678 370927 239699 370957
rect 239678 370923 239694 370927
rect 239870 370923 239886 370957
rect 239954 370929 239975 370957
rect 239954 370923 239970 370929
rect 240146 370923 240162 370957
rect 240230 370929 240251 370957
rect 240230 370923 240246 370929
rect 240422 370923 240438 370957
rect 240506 370931 240527 370957
rect 240506 370923 240522 370931
rect 240698 370923 240714 370957
rect 240782 370929 240803 370957
rect 240782 370923 240798 370929
rect 240974 370923 240990 370957
rect 241058 370929 241079 370957
rect 241058 370923 241074 370929
rect 241250 370923 241266 370957
rect 241334 370929 241357 370957
rect 241334 370923 241350 370929
rect 241526 370923 241542 370957
rect 241610 370929 241633 370957
rect 241610 370923 241626 370929
rect 241802 370923 241818 370957
rect 241886 370927 241905 370957
rect 241886 370923 241902 370927
rect 242078 370923 242094 370957
rect 242162 370927 242183 370957
rect 242162 370923 242178 370927
rect 242354 370923 242370 370957
rect 242438 370931 242459 370957
rect 242438 370923 242454 370931
rect 242630 370923 242646 370957
rect 242714 370933 242737 370957
rect 242714 370923 242730 370933
rect 242906 370923 242922 370957
rect 242990 370929 243011 370957
rect 242990 370923 243006 370929
rect 243182 370923 243198 370957
rect 243266 370933 243287 370957
rect 243266 370923 243282 370933
rect 243458 370923 243474 370957
rect 243542 370933 243565 370957
rect 243542 370923 243558 370933
rect 243734 370923 243750 370957
rect 243818 370935 243841 370957
rect 243818 370923 243834 370935
rect 244010 370923 244026 370957
rect 244094 370931 244117 370957
rect 244094 370923 244110 370931
rect 244286 370923 244302 370957
rect 244370 370933 244393 370957
rect 244370 370923 244386 370933
rect 244562 370923 244578 370957
rect 244646 370933 244669 370957
rect 244646 370923 244662 370933
rect 244838 370923 244854 370957
rect 244922 370935 244943 370957
rect 244922 370923 244938 370935
rect 245114 370923 245130 370957
rect 245198 370935 245223 370957
rect 245198 370923 245214 370935
rect 245390 370923 245406 370957
rect 245474 370935 245499 370957
rect 245474 370923 245490 370935
rect 245666 370923 245682 370957
rect 245750 370935 245771 370957
rect 245750 370923 245766 370935
rect 245942 370923 245958 370957
rect 246026 370925 246047 370957
rect 246026 370923 246042 370925
rect 246218 370923 246234 370957
rect 246302 370923 246318 370957
rect 246494 370923 246510 370957
rect 246578 370925 246609 370957
rect 246740 370999 246774 371015
rect 246578 370923 246594 370925
rect 232648 370873 232682 370889
rect 232648 370797 232682 370813
rect 232806 370873 232840 370889
rect 232806 370797 232840 370813
rect 232924 370873 232958 370889
rect 232924 370797 232958 370813
rect 233082 370873 233116 370889
rect 233082 370797 233116 370813
rect 233200 370873 233234 370889
rect 233200 370797 233234 370813
rect 233358 370873 233392 370889
rect 233358 370797 233392 370813
rect 233476 370873 233510 370889
rect 233476 370797 233510 370813
rect 233634 370873 233668 370889
rect 233634 370797 233668 370813
rect 233752 370873 233786 370889
rect 233752 370797 233786 370813
rect 233910 370873 233944 370889
rect 233910 370797 233944 370813
rect 234028 370873 234062 370889
rect 234028 370797 234062 370813
rect 234186 370873 234220 370889
rect 234186 370797 234220 370813
rect 234304 370873 234338 370889
rect 234304 370797 234338 370813
rect 234462 370873 234496 370889
rect 234462 370797 234496 370813
rect 234580 370873 234614 370889
rect 234580 370797 234614 370813
rect 234738 370873 234772 370889
rect 234738 370797 234772 370813
rect 234856 370873 234890 370889
rect 234856 370797 234890 370813
rect 235014 370873 235048 370889
rect 235014 370797 235048 370813
rect 235132 370873 235166 370889
rect 235132 370797 235166 370813
rect 235290 370873 235324 370889
rect 235290 370797 235324 370813
rect 235408 370873 235442 370889
rect 235408 370797 235442 370813
rect 235566 370873 235600 370889
rect 235566 370797 235600 370813
rect 235684 370873 235718 370889
rect 235684 370797 235718 370813
rect 235842 370873 235876 370889
rect 235842 370797 235876 370813
rect 235960 370873 235994 370889
rect 235960 370797 235994 370813
rect 236118 370873 236152 370889
rect 236118 370797 236152 370813
rect 236236 370873 236270 370889
rect 236236 370797 236270 370813
rect 236394 370873 236428 370889
rect 236394 370797 236428 370813
rect 236512 370873 236546 370889
rect 236512 370797 236546 370813
rect 236670 370873 236704 370889
rect 236670 370797 236704 370813
rect 236788 370873 236822 370889
rect 236788 370797 236822 370813
rect 236946 370873 236980 370889
rect 236946 370797 236980 370813
rect 237064 370873 237098 370889
rect 237064 370797 237098 370813
rect 237222 370873 237256 370889
rect 237222 370797 237256 370813
rect 237340 370873 237374 370889
rect 237340 370797 237374 370813
rect 237498 370873 237532 370889
rect 237498 370797 237532 370813
rect 237616 370873 237650 370889
rect 237616 370797 237650 370813
rect 237774 370873 237808 370889
rect 237774 370797 237808 370813
rect 237892 370873 237926 370889
rect 237892 370797 237926 370813
rect 238050 370873 238084 370889
rect 238050 370797 238084 370813
rect 238168 370873 238202 370889
rect 238168 370797 238202 370813
rect 238326 370873 238360 370889
rect 238326 370797 238360 370813
rect 238444 370873 238478 370889
rect 238444 370797 238478 370813
rect 238602 370873 238636 370889
rect 238602 370797 238636 370813
rect 238720 370873 238754 370889
rect 238720 370797 238754 370813
rect 238878 370873 238912 370889
rect 238878 370797 238912 370813
rect 238996 370873 239030 370889
rect 238996 370797 239030 370813
rect 239154 370873 239188 370889
rect 239154 370797 239188 370813
rect 239272 370873 239306 370889
rect 239272 370797 239306 370813
rect 239430 370873 239464 370889
rect 239430 370797 239464 370813
rect 239548 370873 239582 370889
rect 239548 370797 239582 370813
rect 239706 370873 239740 370889
rect 239706 370797 239740 370813
rect 239824 370873 239858 370889
rect 239824 370797 239858 370813
rect 239982 370873 240016 370889
rect 239982 370797 240016 370813
rect 240100 370873 240134 370889
rect 240100 370797 240134 370813
rect 240258 370873 240292 370889
rect 240258 370797 240292 370813
rect 240376 370873 240410 370889
rect 240376 370797 240410 370813
rect 240534 370873 240568 370889
rect 240534 370797 240568 370813
rect 240652 370873 240686 370889
rect 240652 370797 240686 370813
rect 240810 370873 240844 370889
rect 240810 370797 240844 370813
rect 240928 370873 240962 370889
rect 240928 370797 240962 370813
rect 241086 370873 241120 370889
rect 241086 370797 241120 370813
rect 241204 370873 241238 370889
rect 241204 370797 241238 370813
rect 241362 370873 241396 370889
rect 241362 370797 241396 370813
rect 241480 370873 241514 370889
rect 241480 370797 241514 370813
rect 241638 370873 241672 370889
rect 241638 370797 241672 370813
rect 241756 370873 241790 370889
rect 241756 370797 241790 370813
rect 241914 370873 241948 370889
rect 241914 370797 241948 370813
rect 242032 370873 242066 370889
rect 242032 370797 242066 370813
rect 242190 370873 242224 370889
rect 242190 370797 242224 370813
rect 242308 370873 242342 370889
rect 242308 370797 242342 370813
rect 242466 370873 242500 370889
rect 242466 370797 242500 370813
rect 242584 370873 242618 370889
rect 242584 370797 242618 370813
rect 242742 370873 242776 370889
rect 242742 370797 242776 370813
rect 242860 370873 242894 370889
rect 242860 370797 242894 370813
rect 243018 370873 243052 370889
rect 243018 370797 243052 370813
rect 243136 370873 243170 370889
rect 243136 370797 243170 370813
rect 243294 370873 243328 370889
rect 243294 370797 243328 370813
rect 243412 370873 243446 370889
rect 243412 370797 243446 370813
rect 243570 370873 243604 370889
rect 243570 370797 243604 370813
rect 243688 370873 243722 370889
rect 243688 370797 243722 370813
rect 243846 370873 243880 370889
rect 243846 370797 243880 370813
rect 243964 370873 243998 370889
rect 243964 370797 243998 370813
rect 244122 370873 244156 370889
rect 244122 370797 244156 370813
rect 244240 370873 244274 370889
rect 244240 370797 244274 370813
rect 244398 370873 244432 370889
rect 244398 370797 244432 370813
rect 244516 370873 244550 370889
rect 244516 370797 244550 370813
rect 244674 370873 244708 370889
rect 244674 370797 244708 370813
rect 244792 370873 244826 370889
rect 244792 370797 244826 370813
rect 244950 370873 244984 370889
rect 244950 370797 244984 370813
rect 245068 370873 245102 370889
rect 245068 370797 245102 370813
rect 245226 370873 245260 370889
rect 245226 370797 245260 370813
rect 245344 370873 245378 370889
rect 245344 370797 245378 370813
rect 245502 370873 245536 370889
rect 245502 370797 245536 370813
rect 245620 370873 245654 370889
rect 245620 370797 245654 370813
rect 245778 370873 245812 370889
rect 245778 370797 245812 370813
rect 245896 370873 245930 370889
rect 245896 370797 245930 370813
rect 246054 370873 246088 370889
rect 246054 370797 246088 370813
rect 246172 370873 246206 370889
rect 246172 370797 246206 370813
rect 246330 370873 246364 370889
rect 246330 370797 246364 370813
rect 246448 370873 246482 370889
rect 246448 370797 246482 370813
rect 246606 370873 246640 370889
rect 246606 370797 246640 370813
rect 232694 370729 232710 370763
rect 232778 370760 232794 370763
rect 232778 370729 232802 370760
rect 232970 370729 232986 370763
rect 233054 370729 233070 370763
rect 233246 370759 233262 370763
rect 233243 370729 233262 370759
rect 233330 370729 233346 370763
rect 233522 370755 233538 370763
rect 233519 370729 233538 370755
rect 233606 370729 233622 370763
rect 233798 370749 233814 370763
rect 233797 370729 233814 370749
rect 233882 370729 233898 370763
rect 234074 370745 234090 370763
rect 234073 370729 234090 370745
rect 234158 370729 234174 370763
rect 234350 370747 234366 370763
rect 234347 370729 234366 370747
rect 234434 370729 234450 370763
rect 234626 370745 234642 370763
rect 234625 370729 234642 370745
rect 234710 370729 234726 370763
rect 234902 370729 234918 370763
rect 234986 370729 235002 370763
rect 235178 370745 235194 370763
rect 235177 370729 235194 370745
rect 235262 370729 235278 370763
rect 235454 370729 235470 370763
rect 235538 370729 235554 370763
rect 235730 370755 235746 370763
rect 235727 370739 235746 370755
rect 235726 370729 235746 370739
rect 235814 370729 235830 370763
rect 236006 370755 236022 370763
rect 236003 370729 236022 370755
rect 236090 370729 236106 370763
rect 236282 370729 236298 370763
rect 236366 370729 236382 370763
rect 236558 370749 236574 370763
rect 236551 370729 236574 370749
rect 236642 370729 236658 370763
rect 236834 370729 236850 370763
rect 236918 370729 236934 370763
rect 237110 370749 237126 370763
rect 237109 370729 237126 370749
rect 237194 370729 237210 370763
rect 237386 370745 237402 370763
rect 237385 370729 237402 370745
rect 237470 370729 237486 370763
rect 237662 370753 237678 370763
rect 237659 370729 237678 370753
rect 237746 370729 237762 370763
rect 237938 370745 237954 370763
rect 237937 370729 237954 370745
rect 238022 370729 238038 370763
rect 238214 370747 238230 370763
rect 238207 370729 238230 370747
rect 238298 370729 238314 370763
rect 238490 370753 238506 370763
rect 238483 370729 238506 370753
rect 238574 370729 238590 370763
rect 238766 370759 238782 370763
rect 238765 370729 238782 370759
rect 238850 370729 238866 370763
rect 239042 370755 239058 370763
rect 239041 370729 239058 370755
rect 239126 370729 239142 370763
rect 239318 370755 239334 370763
rect 239315 370729 239334 370755
rect 239402 370729 239418 370763
rect 239594 370755 239610 370763
rect 239587 370729 239610 370755
rect 239678 370729 239694 370763
rect 239870 370755 239886 370763
rect 239869 370729 239886 370755
rect 239954 370729 239970 370763
rect 240146 370729 240162 370763
rect 240230 370729 240246 370763
rect 240422 370749 240438 370763
rect 240421 370729 240438 370749
rect 240506 370729 240522 370763
rect 240698 370729 240714 370763
rect 240782 370729 240798 370763
rect 240974 370729 240990 370763
rect 241058 370729 241074 370763
rect 241250 370741 241266 370763
rect 241243 370729 241266 370741
rect 241334 370729 241350 370763
rect 241526 370737 241542 370763
rect 241525 370729 241542 370737
rect 241610 370729 241626 370763
rect 241802 370729 241818 370763
rect 241886 370729 241902 370763
rect 242078 370737 242094 370763
rect 242077 370729 242094 370737
rect 242162 370729 242178 370763
rect 242354 370737 242370 370763
rect 242353 370729 242370 370737
rect 242438 370729 242454 370763
rect 242630 370753 242646 370763
rect 242623 370729 242646 370753
rect 242714 370729 242730 370763
rect 242906 370745 242922 370763
rect 242901 370729 242922 370745
rect 242990 370729 243006 370763
rect 243182 370729 243198 370763
rect 243266 370729 243282 370763
rect 243458 370729 243474 370763
rect 243542 370745 243558 370763
rect 243734 370749 243750 370763
rect 243542 370729 243563 370745
rect 232700 370520 232802 370729
rect 232971 370520 233069 370729
rect 233243 370520 233341 370729
rect 233519 370520 233617 370729
rect 233797 370520 233895 370729
rect 234073 370520 234171 370729
rect 234347 370520 234445 370729
rect 234625 370520 234723 370729
rect 234903 370520 235001 370729
rect 235177 370520 235275 370729
rect 235455 370520 235553 370729
rect 235726 370520 235826 370729
rect 236003 370520 236101 370729
rect 236283 370520 236381 370729
rect 236551 370520 236649 370729
rect 236835 370520 236933 370729
rect 237109 370520 237207 370729
rect 237385 370520 237483 370729
rect 237659 370520 237757 370729
rect 237937 370520 238035 370729
rect 238207 370520 238305 370729
rect 238483 370520 238581 370729
rect 238765 370520 238863 370729
rect 239041 370520 239139 370729
rect 239315 370714 239413 370729
rect 239587 370520 239685 370729
rect 239869 370520 239967 370729
rect 240147 370520 240245 370729
rect 240421 370520 240519 370729
rect 240699 370520 240797 370729
rect 240975 370520 241073 370729
rect 241243 370520 241341 370729
rect 241525 370520 241623 370729
rect 241803 370520 241901 370729
rect 242077 370520 242175 370729
rect 242353 370520 242451 370729
rect 242623 370520 242721 370729
rect 242901 370520 242999 370729
rect 243183 370520 243281 370729
rect 243465 370520 243563 370729
rect 243733 370729 243750 370749
rect 243818 370729 243834 370763
rect 244010 370749 244026 370763
rect 244009 370729 244026 370749
rect 244094 370729 244110 370763
rect 244286 370749 244302 370763
rect 244279 370729 244302 370749
rect 244370 370729 244386 370763
rect 244562 370755 244578 370763
rect 244557 370729 244578 370755
rect 244646 370729 244662 370763
rect 244838 370729 244854 370763
rect 244922 370729 244938 370763
rect 245114 370729 245130 370763
rect 245198 370755 245214 370763
rect 245198 370729 245217 370755
rect 245390 370753 245406 370763
rect 243733 370520 243831 370729
rect 244009 370520 244107 370729
rect 244279 370520 244377 370729
rect 244557 370520 244655 370729
rect 244839 370520 244937 370729
rect 245119 370520 245217 370729
rect 245385 370729 245406 370753
rect 245474 370729 245490 370763
rect 245666 370747 245682 370763
rect 245661 370729 245682 370747
rect 245750 370729 245766 370763
rect 245942 370753 245958 370763
rect 245941 370729 245958 370753
rect 246026 370729 246042 370763
rect 246218 370729 246234 370763
rect 246302 370753 246318 370763
rect 246302 370729 246323 370753
rect 246494 370729 246510 370763
rect 246578 370757 246594 370763
rect 246578 370729 246601 370757
rect 245385 370520 245483 370729
rect 245661 370520 245759 370729
rect 245941 370520 246039 370729
rect 246225 370520 246323 370729
rect 246503 370520 246601 370729
rect 246740 370671 246774 370687
rect 247092 370520 247190 371144
rect 232697 370489 247190 370520
rect 232697 370433 236703 370489
rect 236781 370433 247190 370489
rect 232697 370422 247190 370433
rect 234266 252206 234346 252216
rect 234266 252164 234282 252206
rect 234336 252164 234346 252206
rect 234266 251839 234346 252164
rect 234539 252096 248751 252123
rect 234538 252025 248751 252096
rect 234538 251839 234636 252025
rect 234814 251839 234912 252025
rect 235088 251839 235186 252025
rect 235366 251839 235464 252025
rect 235638 251839 235736 252025
rect 235916 251839 236014 252025
rect 236194 251839 236292 252025
rect 236472 251839 236570 252025
rect 236746 251839 236844 252025
rect 237022 251839 237120 252025
rect 237298 251839 237396 252025
rect 237576 251839 237674 252025
rect 237852 251839 237950 252025
rect 238124 251839 238222 252025
rect 238402 251839 238500 252025
rect 238674 251839 238772 252025
rect 238952 251839 239050 252025
rect 239228 251839 239326 252025
rect 234255 251805 234271 251839
rect 234339 251805 234355 251839
rect 234531 251805 234547 251839
rect 234615 251814 234636 251839
rect 234615 251805 234631 251814
rect 234807 251805 234823 251839
rect 234891 251816 234912 251839
rect 234891 251805 234907 251816
rect 235083 251805 235099 251839
rect 235167 251812 235186 251839
rect 235167 251805 235183 251812
rect 235359 251805 235375 251839
rect 235443 251812 235464 251839
rect 235443 251805 235459 251812
rect 235635 251805 235651 251839
rect 235719 251814 235736 251839
rect 235719 251805 235735 251814
rect 235911 251805 235927 251839
rect 235995 251812 236014 251839
rect 235995 251805 236011 251812
rect 236187 251805 236203 251839
rect 236271 251812 236292 251839
rect 236271 251805 236287 251812
rect 236463 251805 236479 251839
rect 236547 251816 236570 251839
rect 236547 251805 236563 251816
rect 236739 251805 236755 251839
rect 236823 251812 236844 251839
rect 236823 251805 236839 251812
rect 237015 251805 237031 251839
rect 237099 251816 237120 251839
rect 237099 251805 237115 251816
rect 237291 251805 237307 251839
rect 237375 251816 237396 251839
rect 237375 251805 237391 251816
rect 237567 251805 237583 251839
rect 237651 251818 237674 251839
rect 237651 251805 237667 251818
rect 237843 251805 237859 251839
rect 237927 251808 237950 251839
rect 237927 251805 237943 251808
rect 238119 251805 238135 251839
rect 238203 251812 238222 251839
rect 238203 251805 238219 251812
rect 238395 251805 238411 251839
rect 238479 251812 238500 251839
rect 238479 251805 238495 251812
rect 238671 251805 238687 251839
rect 238755 251805 238772 251839
rect 238947 251805 238963 251839
rect 239031 251812 239050 251839
rect 239031 251805 239047 251812
rect 239223 251805 239239 251839
rect 239307 251812 239326 251839
rect 239498 251839 239596 252025
rect 239784 251839 239882 252025
rect 240056 251839 240154 252025
rect 240336 251839 240434 252025
rect 240610 251839 240708 252025
rect 240886 251839 240984 252025
rect 241162 251839 241260 252025
rect 241438 251839 241536 252025
rect 241714 251839 241812 252025
rect 241990 251839 242088 252025
rect 242266 251839 242364 252025
rect 242542 251839 242640 252025
rect 242820 251839 242918 252025
rect 243096 251839 243194 252025
rect 243368 251839 243466 252025
rect 243646 251839 243744 252025
rect 243922 251839 244020 252025
rect 244200 251839 244298 252025
rect 244474 251839 244572 252025
rect 244750 251839 244848 252025
rect 245028 251839 245126 252025
rect 245304 251839 245402 252025
rect 245580 251839 245678 252025
rect 245856 251839 245954 252025
rect 246132 251839 246230 252025
rect 246406 251839 246504 252025
rect 246686 251839 246784 252025
rect 246962 251839 247060 252025
rect 247234 251839 247332 252025
rect 247510 251839 247608 252025
rect 247780 251839 247878 252025
rect 248072 251839 248170 252025
rect 239307 251805 239323 251812
rect 239498 251810 239515 251839
rect 239499 251805 239515 251810
rect 239583 251805 239599 251839
rect 239775 251805 239791 251839
rect 239859 251808 239882 251839
rect 239859 251805 239875 251808
rect 240051 251805 240067 251839
rect 240135 251808 240154 251839
rect 240135 251805 240151 251808
rect 240327 251805 240343 251839
rect 240411 251808 240434 251839
rect 240411 251805 240427 251808
rect 240603 251805 240619 251839
rect 240687 251808 240708 251839
rect 240687 251805 240703 251808
rect 240879 251805 240895 251839
rect 240963 251810 240984 251839
rect 240963 251805 240979 251810
rect 241155 251805 241171 251839
rect 241239 251808 241260 251839
rect 241239 251805 241255 251808
rect 241431 251805 241447 251839
rect 241515 251810 241536 251839
rect 241515 251805 241531 251810
rect 241707 251805 241723 251839
rect 241791 251810 241812 251839
rect 241791 251805 241807 251810
rect 241983 251805 241999 251839
rect 242067 251812 242088 251839
rect 242067 251805 242083 251812
rect 242259 251805 242275 251839
rect 242343 251810 242364 251839
rect 242343 251805 242359 251810
rect 242535 251805 242551 251839
rect 242619 251810 242640 251839
rect 242619 251805 242635 251810
rect 242811 251805 242827 251839
rect 242895 251810 242918 251839
rect 242895 251805 242911 251810
rect 243087 251805 243103 251839
rect 243171 251810 243194 251839
rect 243171 251805 243187 251810
rect 243363 251805 243379 251839
rect 243447 251808 243466 251839
rect 243447 251805 243463 251808
rect 243639 251805 243655 251839
rect 243723 251808 243744 251839
rect 243723 251805 243739 251808
rect 243915 251805 243931 251839
rect 243999 251812 244020 251839
rect 243999 251805 244015 251812
rect 244191 251805 244207 251839
rect 244275 251814 244298 251839
rect 244275 251805 244291 251814
rect 244467 251805 244483 251839
rect 244551 251810 244572 251839
rect 244551 251805 244567 251810
rect 244743 251805 244759 251839
rect 244827 251814 244848 251839
rect 244827 251805 244843 251814
rect 245019 251805 245035 251839
rect 245103 251814 245126 251839
rect 245103 251805 245119 251814
rect 245295 251805 245311 251839
rect 245379 251816 245402 251839
rect 245379 251805 245395 251816
rect 245571 251805 245587 251839
rect 245655 251812 245678 251839
rect 245655 251805 245671 251812
rect 245847 251805 245863 251839
rect 245931 251814 245954 251839
rect 245931 251805 245947 251814
rect 246123 251805 246139 251839
rect 246207 251814 246230 251839
rect 246207 251805 246223 251814
rect 246399 251805 246415 251839
rect 246483 251816 246504 251839
rect 246483 251805 246499 251816
rect 246675 251805 246691 251839
rect 246759 251816 246784 251839
rect 246759 251805 246775 251816
rect 246951 251805 246967 251839
rect 247035 251816 247060 251839
rect 247035 251805 247051 251816
rect 247227 251805 247243 251839
rect 247311 251816 247332 251839
rect 247311 251805 247327 251816
rect 247503 251805 247519 251839
rect 247587 251806 247608 251839
rect 247587 251805 247603 251806
rect 247779 251805 247795 251839
rect 247863 251805 247879 251839
rect 248055 251805 248071 251839
rect 248139 251806 248170 251839
rect 248301 251881 248335 251897
rect 248139 251805 248155 251806
rect 234266 251800 234346 251805
rect 238674 251804 238772 251805
rect 247780 251804 247878 251805
rect 147704 251784 150583 251795
rect 147704 251753 150584 251784
rect 58707 251582 60075 251618
rect 58707 251246 58743 251582
rect 58907 251515 58977 251582
rect 59175 251515 59245 251582
rect 59723 251515 59793 251582
rect 60005 251515 60075 251582
rect 60236 251557 60270 251573
rect 58886 251481 58902 251515
rect 58970 251481 58986 251515
rect 59162 251481 59178 251515
rect 59246 251481 59262 251515
rect 59438 251481 59454 251515
rect 59522 251481 59538 251515
rect 59714 251481 59730 251515
rect 59798 251481 59814 251515
rect 59990 251481 60006 251515
rect 60074 251481 60090 251515
rect 58907 251476 58977 251481
rect 59175 251476 59245 251481
rect 59723 251474 59793 251481
rect 60005 251476 60075 251481
rect 58840 251431 58874 251447
rect 58840 251355 58874 251371
rect 58998 251431 59032 251447
rect 58998 251355 59032 251371
rect 59116 251431 59150 251447
rect 59116 251355 59150 251371
rect 59274 251431 59308 251447
rect 59274 251355 59308 251371
rect 59392 251431 59426 251447
rect 59392 251355 59426 251371
rect 59550 251431 59584 251447
rect 59550 251355 59584 251371
rect 59668 251431 59702 251447
rect 59668 251355 59702 251371
rect 59826 251431 59860 251447
rect 59826 251355 59860 251371
rect 59944 251431 59978 251447
rect 59944 251355 59978 251371
rect 60102 251431 60136 251447
rect 60102 251355 60136 251371
rect 59721 251321 59817 251322
rect 58886 251287 58902 251321
rect 58970 251287 58986 251321
rect 59162 251287 59178 251321
rect 59246 251287 59262 251321
rect 59438 251287 59454 251321
rect 59522 251287 59538 251321
rect 59714 251287 59730 251321
rect 59798 251287 59817 251321
rect 59990 251287 60006 251321
rect 60074 251287 60090 251321
rect 59165 251246 59259 251287
rect 59721 251250 59817 251287
rect 60011 251260 60075 251287
rect 60011 251250 60073 251260
rect 59719 251246 60073 251250
rect 58707 251244 60073 251246
rect 58707 251210 58923 251244
rect 58961 251210 60073 251244
rect 147704 251310 147746 251753
rect 148024 251748 150584 251753
rect 148024 251639 148102 251748
rect 148300 251639 148378 251748
rect 148578 251639 148656 251748
rect 148850 251639 148928 251748
rect 149132 251639 149210 251646
rect 149404 251639 149482 251748
rect 149680 251639 149758 251748
rect 149954 251639 150032 251748
rect 150232 251639 150310 251748
rect 150506 251639 150584 251748
rect 234209 251755 234243 251771
rect 150741 251681 150775 251697
rect 148011 251605 148027 251639
rect 148095 251605 148111 251639
rect 148287 251605 148303 251639
rect 148371 251605 148387 251639
rect 148563 251605 148579 251639
rect 148647 251605 148663 251639
rect 148839 251605 148855 251639
rect 148923 251605 148939 251639
rect 149115 251605 149131 251639
rect 149199 251605 149215 251639
rect 149391 251605 149407 251639
rect 149475 251605 149491 251639
rect 149667 251605 149683 251639
rect 149751 251605 149767 251639
rect 149943 251605 149959 251639
rect 150027 251605 150043 251639
rect 150219 251605 150235 251639
rect 150303 251605 150319 251639
rect 150495 251605 150511 251639
rect 150579 251605 150595 251639
rect 148024 251604 148102 251605
rect 148300 251602 148378 251605
rect 148578 251604 148656 251605
rect 148850 251604 148928 251605
rect 149132 251604 149210 251605
rect 149404 251604 149482 251605
rect 149680 251602 149758 251605
rect 149954 251602 150032 251605
rect 150232 251604 150310 251605
rect 150506 251602 150584 251605
rect 147965 251555 147999 251571
rect 147965 251479 147999 251495
rect 148123 251555 148157 251571
rect 148123 251479 148157 251495
rect 148241 251555 148275 251571
rect 148241 251479 148275 251495
rect 148399 251555 148433 251571
rect 148399 251479 148433 251495
rect 148517 251555 148551 251571
rect 148517 251479 148551 251495
rect 148675 251555 148709 251571
rect 148675 251479 148709 251495
rect 148793 251555 148827 251571
rect 148793 251479 148827 251495
rect 148951 251555 148985 251571
rect 148951 251479 148985 251495
rect 149069 251555 149103 251571
rect 149069 251479 149103 251495
rect 149227 251555 149261 251571
rect 149227 251479 149261 251495
rect 149345 251555 149379 251571
rect 149345 251479 149379 251495
rect 149503 251555 149537 251571
rect 149503 251479 149537 251495
rect 149621 251555 149655 251571
rect 149621 251479 149655 251495
rect 149779 251555 149813 251571
rect 149779 251479 149813 251495
rect 149897 251555 149931 251571
rect 149897 251479 149931 251495
rect 150055 251555 150089 251571
rect 150055 251479 150089 251495
rect 150173 251555 150207 251571
rect 150173 251479 150207 251495
rect 150331 251555 150365 251571
rect 150331 251479 150365 251495
rect 150449 251555 150483 251571
rect 150449 251479 150483 251495
rect 150607 251555 150641 251571
rect 150607 251479 150641 251495
rect 148028 251445 148106 251446
rect 148854 251445 148932 251446
rect 149130 251445 149208 251446
rect 149402 251445 149480 251448
rect 149680 251445 149758 251446
rect 149958 251445 150036 251448
rect 150234 251445 150312 251448
rect 150510 251445 150588 251450
rect 148011 251411 148027 251445
rect 148095 251411 148111 251445
rect 148287 251411 148303 251445
rect 148371 251411 148387 251445
rect 148563 251411 148579 251445
rect 148647 251411 148663 251445
rect 148839 251411 148855 251445
rect 148923 251411 148939 251445
rect 149115 251411 149131 251445
rect 149199 251411 149215 251445
rect 149391 251411 149407 251445
rect 149475 251411 149491 251445
rect 149667 251411 149683 251445
rect 149751 251411 149767 251445
rect 149943 251411 149959 251445
rect 150027 251411 150043 251445
rect 150219 251411 150235 251445
rect 150303 251411 150319 251445
rect 150495 251411 150511 251445
rect 150579 251411 150595 251445
rect 148028 251310 148106 251411
rect 148302 251310 148380 251411
rect 148578 251310 148656 251411
rect 148854 251310 148932 251411
rect 149130 251404 149208 251411
rect 149402 251310 149480 251411
rect 149680 251310 149758 251411
rect 149958 251310 150036 251411
rect 150234 251310 150312 251411
rect 150510 251310 150588 251411
rect 234209 251679 234243 251695
rect 234367 251755 234401 251771
rect 234367 251679 234401 251695
rect 234485 251755 234519 251771
rect 234485 251679 234519 251695
rect 234643 251755 234677 251771
rect 234643 251679 234677 251695
rect 234761 251755 234795 251771
rect 234761 251679 234795 251695
rect 234919 251755 234953 251771
rect 234919 251679 234953 251695
rect 235037 251755 235071 251771
rect 235037 251679 235071 251695
rect 235195 251755 235229 251771
rect 235195 251679 235229 251695
rect 235313 251755 235347 251771
rect 235313 251679 235347 251695
rect 235471 251755 235505 251771
rect 235471 251679 235505 251695
rect 235589 251755 235623 251771
rect 235589 251679 235623 251695
rect 235747 251755 235781 251771
rect 235747 251679 235781 251695
rect 235865 251755 235899 251771
rect 235865 251679 235899 251695
rect 236023 251755 236057 251771
rect 236023 251679 236057 251695
rect 236141 251755 236175 251771
rect 236141 251679 236175 251695
rect 236299 251755 236333 251771
rect 236299 251679 236333 251695
rect 236417 251755 236451 251771
rect 236417 251679 236451 251695
rect 236575 251755 236609 251771
rect 236575 251679 236609 251695
rect 236693 251755 236727 251771
rect 236693 251679 236727 251695
rect 236851 251755 236885 251771
rect 236851 251679 236885 251695
rect 236969 251755 237003 251771
rect 236969 251679 237003 251695
rect 237127 251755 237161 251771
rect 237127 251679 237161 251695
rect 237245 251755 237279 251771
rect 237245 251679 237279 251695
rect 237403 251755 237437 251771
rect 237403 251679 237437 251695
rect 237521 251755 237555 251771
rect 237521 251679 237555 251695
rect 237679 251755 237713 251771
rect 237679 251679 237713 251695
rect 237797 251755 237831 251771
rect 237797 251679 237831 251695
rect 237955 251755 237989 251771
rect 237955 251679 237989 251695
rect 238073 251755 238107 251771
rect 238073 251679 238107 251695
rect 238231 251755 238265 251771
rect 238231 251679 238265 251695
rect 238349 251755 238383 251771
rect 238349 251679 238383 251695
rect 238507 251755 238541 251771
rect 238507 251679 238541 251695
rect 238625 251755 238659 251771
rect 238625 251679 238659 251695
rect 238783 251755 238817 251771
rect 238783 251679 238817 251695
rect 238901 251755 238935 251771
rect 238901 251679 238935 251695
rect 239059 251755 239093 251771
rect 239059 251679 239093 251695
rect 239177 251755 239211 251771
rect 239177 251679 239211 251695
rect 239335 251755 239369 251771
rect 239335 251679 239369 251695
rect 239453 251755 239487 251771
rect 239453 251679 239487 251695
rect 239611 251755 239645 251771
rect 239611 251679 239645 251695
rect 239729 251755 239763 251771
rect 239729 251679 239763 251695
rect 239887 251755 239921 251771
rect 239887 251679 239921 251695
rect 240005 251755 240039 251771
rect 240005 251679 240039 251695
rect 240163 251755 240197 251771
rect 240163 251679 240197 251695
rect 240281 251755 240315 251771
rect 240281 251679 240315 251695
rect 240439 251755 240473 251771
rect 240439 251679 240473 251695
rect 240557 251755 240591 251771
rect 240557 251679 240591 251695
rect 240715 251755 240749 251771
rect 240715 251679 240749 251695
rect 240833 251755 240867 251771
rect 240833 251679 240867 251695
rect 240991 251755 241025 251771
rect 240991 251679 241025 251695
rect 241109 251755 241143 251771
rect 241109 251679 241143 251695
rect 241267 251755 241301 251771
rect 241267 251679 241301 251695
rect 241385 251755 241419 251771
rect 241385 251679 241419 251695
rect 241543 251755 241577 251771
rect 241543 251679 241577 251695
rect 241661 251755 241695 251771
rect 241661 251679 241695 251695
rect 241819 251755 241853 251771
rect 241819 251679 241853 251695
rect 241937 251755 241971 251771
rect 241937 251679 241971 251695
rect 242095 251755 242129 251771
rect 242095 251679 242129 251695
rect 242213 251755 242247 251771
rect 242213 251679 242247 251695
rect 242371 251755 242405 251771
rect 242371 251679 242405 251695
rect 242489 251755 242523 251771
rect 242489 251679 242523 251695
rect 242647 251755 242681 251771
rect 242647 251679 242681 251695
rect 242765 251755 242799 251771
rect 242765 251679 242799 251695
rect 242923 251755 242957 251771
rect 242923 251679 242957 251695
rect 243041 251755 243075 251771
rect 243041 251679 243075 251695
rect 243199 251755 243233 251771
rect 243199 251679 243233 251695
rect 243317 251755 243351 251771
rect 243317 251679 243351 251695
rect 243475 251755 243509 251771
rect 243475 251679 243509 251695
rect 243593 251755 243627 251771
rect 243593 251679 243627 251695
rect 243751 251755 243785 251771
rect 243751 251679 243785 251695
rect 243869 251755 243903 251771
rect 243869 251679 243903 251695
rect 244027 251755 244061 251771
rect 244027 251679 244061 251695
rect 244145 251755 244179 251771
rect 244145 251679 244179 251695
rect 244303 251755 244337 251771
rect 244303 251679 244337 251695
rect 244421 251755 244455 251771
rect 244421 251679 244455 251695
rect 244579 251755 244613 251771
rect 244579 251679 244613 251695
rect 244697 251755 244731 251771
rect 244697 251679 244731 251695
rect 244855 251755 244889 251771
rect 244855 251679 244889 251695
rect 244973 251755 245007 251771
rect 244973 251679 245007 251695
rect 245131 251755 245165 251771
rect 245131 251679 245165 251695
rect 245249 251755 245283 251771
rect 245249 251679 245283 251695
rect 245407 251755 245441 251771
rect 245407 251679 245441 251695
rect 245525 251755 245559 251771
rect 245525 251679 245559 251695
rect 245683 251755 245717 251771
rect 245683 251679 245717 251695
rect 245801 251755 245835 251771
rect 245801 251679 245835 251695
rect 245959 251755 245993 251771
rect 245959 251679 245993 251695
rect 246077 251755 246111 251771
rect 246077 251679 246111 251695
rect 246235 251755 246269 251771
rect 246235 251679 246269 251695
rect 246353 251755 246387 251771
rect 246353 251679 246387 251695
rect 246511 251755 246545 251771
rect 246511 251679 246545 251695
rect 246629 251755 246663 251771
rect 246629 251679 246663 251695
rect 246787 251755 246821 251771
rect 246787 251679 246821 251695
rect 246905 251755 246939 251771
rect 246905 251679 246939 251695
rect 247063 251755 247097 251771
rect 247063 251679 247097 251695
rect 247181 251755 247215 251771
rect 247181 251679 247215 251695
rect 247339 251755 247373 251771
rect 247339 251679 247373 251695
rect 247457 251755 247491 251771
rect 247457 251679 247491 251695
rect 247615 251755 247649 251771
rect 247615 251679 247649 251695
rect 247733 251755 247767 251771
rect 247733 251679 247767 251695
rect 247891 251755 247925 251771
rect 247891 251679 247925 251695
rect 248009 251755 248043 251771
rect 248009 251679 248043 251695
rect 248167 251755 248201 251771
rect 248167 251679 248201 251695
rect 234266 251645 234346 251648
rect 234255 251611 234271 251645
rect 234339 251611 234355 251645
rect 234531 251611 234547 251645
rect 234615 251611 234631 251645
rect 234807 251640 234823 251645
rect 234804 251611 234823 251640
rect 234891 251611 234907 251645
rect 235083 251636 235099 251645
rect 235080 251611 235099 251636
rect 235167 251611 235183 251645
rect 235359 251630 235375 251645
rect 235358 251611 235375 251630
rect 235443 251611 235459 251645
rect 235635 251626 235651 251645
rect 235634 251611 235651 251626
rect 235719 251611 235735 251645
rect 235911 251628 235927 251645
rect 235908 251611 235927 251628
rect 235995 251611 236011 251645
rect 236187 251626 236203 251645
rect 236186 251611 236203 251626
rect 236271 251611 236287 251645
rect 236463 251611 236479 251645
rect 236547 251611 236563 251645
rect 236739 251626 236755 251645
rect 236738 251611 236755 251626
rect 236823 251611 236839 251645
rect 237015 251611 237031 251645
rect 237099 251611 237115 251645
rect 237291 251636 237307 251645
rect 237288 251611 237307 251636
rect 237375 251611 237391 251645
rect 237567 251636 237583 251645
rect 237564 251611 237583 251636
rect 237651 251611 237667 251645
rect 237843 251611 237859 251645
rect 237927 251611 237943 251645
rect 238119 251630 238135 251645
rect 238112 251611 238135 251630
rect 238203 251611 238219 251645
rect 238395 251611 238411 251645
rect 238479 251611 238495 251645
rect 238671 251630 238687 251645
rect 238670 251611 238687 251630
rect 238755 251611 238771 251645
rect 238947 251626 238963 251645
rect 238946 251611 238963 251626
rect 239031 251611 239047 251645
rect 239223 251634 239239 251645
rect 239220 251611 239239 251634
rect 239307 251611 239323 251645
rect 239499 251626 239515 251645
rect 239498 251611 239515 251626
rect 239583 251611 239599 251645
rect 239775 251628 239791 251645
rect 239768 251611 239791 251628
rect 239859 251611 239875 251645
rect 240051 251634 240067 251645
rect 240044 251611 240067 251634
rect 240135 251611 240151 251645
rect 240327 251640 240343 251645
rect 240326 251611 240343 251640
rect 240411 251611 240427 251645
rect 240603 251636 240619 251645
rect 240602 251611 240619 251636
rect 240687 251611 240703 251645
rect 240879 251636 240895 251645
rect 240876 251611 240895 251636
rect 240963 251611 240979 251645
rect 241155 251636 241171 251645
rect 241148 251611 241171 251636
rect 241239 251611 241255 251645
rect 241431 251636 241447 251645
rect 241430 251611 241447 251636
rect 241515 251611 241531 251645
rect 241707 251611 241723 251645
rect 241791 251611 241807 251645
rect 241983 251630 241999 251645
rect 241982 251611 241999 251630
rect 242067 251611 242083 251645
rect 242259 251611 242275 251645
rect 242343 251611 242359 251645
rect 242535 251611 242551 251645
rect 242619 251611 242635 251645
rect 242811 251622 242827 251645
rect 242804 251611 242827 251622
rect 242895 251611 242911 251645
rect 243087 251618 243103 251645
rect 243086 251611 243103 251618
rect 243171 251611 243187 251645
rect 243363 251611 243379 251645
rect 243447 251611 243463 251645
rect 243639 251618 243655 251645
rect 243638 251611 243655 251618
rect 243723 251611 243739 251645
rect 243915 251618 243931 251645
rect 243914 251611 243931 251618
rect 243999 251611 244015 251645
rect 244191 251634 244207 251645
rect 244184 251611 244207 251634
rect 244275 251611 244291 251645
rect 244467 251626 244483 251645
rect 244462 251611 244483 251626
rect 244551 251611 244567 251645
rect 244743 251611 244759 251645
rect 244827 251611 244843 251645
rect 245019 251611 245035 251645
rect 245103 251626 245119 251645
rect 245295 251630 245311 251645
rect 245103 251611 245124 251626
rect 150741 251353 150775 251369
rect 147704 251268 150590 251310
rect 234266 251294 234346 251611
rect 234532 251401 234630 251611
rect 234804 251401 234902 251611
rect 235080 251401 235178 251611
rect 235358 251401 235456 251611
rect 235634 251401 235732 251611
rect 235908 251401 236006 251611
rect 236186 251401 236284 251611
rect 236464 251401 236562 251611
rect 236738 251401 236836 251611
rect 237016 251401 237114 251611
rect 237288 251401 237386 251611
rect 237564 251401 237662 251611
rect 237844 251401 237942 251611
rect 238112 251401 238210 251611
rect 238396 251401 238494 251611
rect 238670 251401 238768 251611
rect 238946 251401 239044 251611
rect 239220 251401 239318 251611
rect 239498 251401 239596 251611
rect 239768 251401 239866 251611
rect 240044 251401 240142 251611
rect 240326 251401 240424 251611
rect 240602 251401 240700 251611
rect 240876 251401 240974 251611
rect 241148 251401 241246 251611
rect 241430 251401 241528 251611
rect 241708 251401 241806 251611
rect 241982 251401 242080 251611
rect 242260 251401 242358 251611
rect 242536 251401 242634 251611
rect 242804 251401 242902 251611
rect 243086 251401 243184 251611
rect 243364 251401 243462 251611
rect 243638 251401 243736 251611
rect 243914 251401 244012 251611
rect 244184 251401 244282 251611
rect 244462 251401 244560 251611
rect 244744 251401 244842 251611
rect 245026 251401 245124 251611
rect 245294 251611 245311 251630
rect 245379 251611 245395 251645
rect 245571 251630 245587 251645
rect 245570 251611 245587 251630
rect 245655 251611 245671 251645
rect 245847 251630 245863 251645
rect 245840 251611 245863 251630
rect 245931 251611 245947 251645
rect 246123 251636 246139 251645
rect 246118 251611 246139 251636
rect 246207 251611 246223 251645
rect 246399 251611 246415 251645
rect 246483 251611 246499 251645
rect 246675 251611 246691 251645
rect 246759 251636 246775 251645
rect 246759 251611 246778 251636
rect 246951 251634 246967 251645
rect 245294 251401 245392 251611
rect 245570 251401 245668 251611
rect 245840 251401 245938 251611
rect 246118 251401 246216 251611
rect 246400 251401 246498 251611
rect 246680 251401 246778 251611
rect 246946 251611 246967 251634
rect 247035 251611 247051 251645
rect 247227 251628 247243 251645
rect 247222 251611 247243 251628
rect 247311 251611 247327 251645
rect 247503 251634 247519 251645
rect 247502 251611 247519 251634
rect 247587 251611 247603 251645
rect 247779 251611 247795 251645
rect 247863 251634 247879 251645
rect 247863 251611 247884 251634
rect 248055 251611 248071 251645
rect 248139 251638 248155 251645
rect 248139 251611 248162 251638
rect 246946 251401 247044 251611
rect 247222 251401 247320 251611
rect 247502 251401 247600 251611
rect 247786 251401 247884 251611
rect 248064 251401 248162 251611
rect 248301 251553 248335 251569
rect 248653 251401 248751 252025
rect 413336 251780 427833 251838
rect 503336 251780 517833 251838
rect 413335 251740 427833 251780
rect 413335 251553 413422 251740
rect 413620 251553 413718 251740
rect 413896 251553 413994 251740
rect 414170 251553 414268 251740
rect 414448 251553 414546 251740
rect 414720 251553 414818 251740
rect 414998 251553 415096 251740
rect 415276 251553 415374 251740
rect 415554 251553 415652 251740
rect 415828 251553 415926 251740
rect 416104 251553 416202 251740
rect 416389 251553 416484 251740
rect 416658 251553 416756 251740
rect 416934 251553 417032 251740
rect 417206 251553 417304 251740
rect 417484 251553 417582 251740
rect 417756 251553 417854 251740
rect 418034 251553 418132 251740
rect 418310 251553 418408 251740
rect 413335 251530 413353 251553
rect 413337 251519 413353 251530
rect 413421 251519 413437 251553
rect 413613 251519 413629 251553
rect 413697 251529 413718 251553
rect 413697 251519 413713 251529
rect 413889 251519 413905 251553
rect 413973 251531 413994 251553
rect 413973 251519 413989 251531
rect 414165 251519 414181 251553
rect 414249 251527 414268 251553
rect 414249 251519 414265 251527
rect 414441 251519 414457 251553
rect 414525 251527 414546 251553
rect 414525 251519 414541 251527
rect 414717 251519 414733 251553
rect 414801 251529 414818 251553
rect 414801 251519 414817 251529
rect 414993 251519 415009 251553
rect 415077 251527 415096 251553
rect 415077 251519 415093 251527
rect 415269 251519 415285 251553
rect 415353 251527 415374 251553
rect 415353 251519 415369 251527
rect 415545 251519 415561 251553
rect 415629 251531 415652 251553
rect 415629 251519 415645 251531
rect 415821 251519 415837 251553
rect 415905 251527 415926 251553
rect 415905 251519 415921 251527
rect 416097 251519 416113 251553
rect 416181 251531 416202 251553
rect 416181 251519 416197 251531
rect 416373 251519 416389 251553
rect 416457 251530 416484 251553
rect 416457 251519 416473 251530
rect 416649 251519 416665 251553
rect 416733 251533 416756 251553
rect 416733 251519 416749 251533
rect 416925 251519 416941 251553
rect 417009 251523 417032 251553
rect 417009 251519 417025 251523
rect 417201 251519 417217 251553
rect 417285 251527 417304 251553
rect 417285 251519 417301 251527
rect 417477 251519 417493 251553
rect 417561 251527 417582 251553
rect 417561 251519 417577 251527
rect 417753 251519 417769 251553
rect 417837 251519 417854 251553
rect 418029 251519 418045 251553
rect 418113 251527 418132 251553
rect 418113 251519 418129 251527
rect 418305 251519 418321 251553
rect 418389 251527 418408 251553
rect 418580 251553 418678 251740
rect 418866 251553 418964 251740
rect 419138 251553 419236 251740
rect 419418 251553 419516 251740
rect 419692 251553 419790 251740
rect 420244 251553 420342 251740
rect 420520 251553 420618 251740
rect 420796 251553 420894 251740
rect 421072 251553 421170 251740
rect 421348 251553 421446 251740
rect 421624 251553 421722 251740
rect 421902 251553 422000 251740
rect 422178 251553 422276 251740
rect 422450 251553 422548 251740
rect 422728 251553 422826 251740
rect 423004 251553 423102 251740
rect 423282 251553 423380 251740
rect 423556 251553 423654 251740
rect 423832 251553 423930 251740
rect 424110 251553 424208 251740
rect 424386 251553 424484 251740
rect 424662 251553 424760 251740
rect 424938 251553 425036 251740
rect 425214 251553 425312 251740
rect 425488 251553 425586 251740
rect 425768 251553 425866 251740
rect 426044 251553 426142 251740
rect 426316 251553 426414 251740
rect 426592 251553 426690 251740
rect 426862 251553 426960 251740
rect 427154 251553 427252 251740
rect 418389 251519 418405 251527
rect 418580 251525 418597 251553
rect 418581 251519 418597 251525
rect 418665 251519 418681 251553
rect 418857 251519 418873 251553
rect 418941 251523 418964 251553
rect 418941 251519 418957 251523
rect 419133 251519 419149 251553
rect 419217 251523 419236 251553
rect 419217 251519 419233 251523
rect 419409 251519 419425 251553
rect 419493 251523 419516 251553
rect 419493 251519 419509 251523
rect 419685 251519 419701 251553
rect 419769 251523 419790 251553
rect 419769 251519 419785 251523
rect 419961 251519 419977 251553
rect 420045 251519 420061 251553
rect 420237 251519 420253 251553
rect 420321 251523 420342 251553
rect 420321 251519 420337 251523
rect 420513 251519 420529 251553
rect 420597 251525 420618 251553
rect 420597 251519 420613 251525
rect 420789 251519 420805 251553
rect 420873 251525 420894 251553
rect 420873 251519 420889 251525
rect 421065 251519 421081 251553
rect 421149 251527 421170 251553
rect 421149 251519 421165 251527
rect 421341 251519 421357 251553
rect 421425 251525 421446 251553
rect 421425 251519 421441 251525
rect 421617 251519 421633 251553
rect 421701 251525 421722 251553
rect 421701 251519 421717 251525
rect 421893 251519 421909 251553
rect 421977 251525 422000 251553
rect 421977 251519 421993 251525
rect 422169 251519 422185 251553
rect 422253 251525 422276 251553
rect 422253 251519 422269 251525
rect 422445 251519 422461 251553
rect 422529 251523 422548 251553
rect 422529 251519 422545 251523
rect 422721 251519 422737 251553
rect 422805 251523 422826 251553
rect 422805 251519 422821 251523
rect 422997 251519 423013 251553
rect 423081 251527 423102 251553
rect 423081 251519 423097 251527
rect 423273 251519 423289 251553
rect 423357 251529 423380 251553
rect 423357 251519 423373 251529
rect 423549 251519 423565 251553
rect 423633 251525 423654 251553
rect 423633 251519 423649 251525
rect 423825 251519 423841 251553
rect 423909 251529 423930 251553
rect 423909 251519 423925 251529
rect 424101 251519 424117 251553
rect 424185 251529 424208 251553
rect 424185 251519 424201 251529
rect 424377 251519 424393 251553
rect 424461 251531 424484 251553
rect 424461 251519 424477 251531
rect 424653 251519 424669 251553
rect 424737 251527 424760 251553
rect 424737 251519 424753 251527
rect 424929 251519 424945 251553
rect 425013 251529 425036 251553
rect 425013 251519 425029 251529
rect 425205 251519 425221 251553
rect 425289 251529 425312 251553
rect 425289 251519 425305 251529
rect 425481 251519 425497 251553
rect 425565 251531 425586 251553
rect 425565 251519 425581 251531
rect 425757 251519 425773 251553
rect 425841 251531 425866 251553
rect 425841 251519 425857 251531
rect 426033 251519 426049 251553
rect 426117 251531 426142 251553
rect 426117 251519 426133 251531
rect 426309 251519 426325 251553
rect 426393 251531 426414 251553
rect 426393 251519 426409 251531
rect 426585 251519 426601 251553
rect 426669 251521 426690 251553
rect 426669 251519 426685 251521
rect 426861 251519 426877 251553
rect 426945 251519 426961 251553
rect 427137 251519 427153 251553
rect 427221 251521 427252 251553
rect 427383 251595 427417 251611
rect 427221 251519 427237 251521
rect 234532 251370 248751 251401
rect 413291 251469 413325 251485
rect 413291 251393 413325 251409
rect 413449 251469 413483 251485
rect 413449 251393 413483 251409
rect 413567 251469 413601 251485
rect 413567 251393 413601 251409
rect 413725 251469 413759 251485
rect 413725 251393 413759 251409
rect 413843 251469 413877 251485
rect 413843 251393 413877 251409
rect 414001 251469 414035 251485
rect 414001 251393 414035 251409
rect 414119 251469 414153 251485
rect 414119 251393 414153 251409
rect 414277 251469 414311 251485
rect 414277 251393 414311 251409
rect 414395 251469 414429 251485
rect 414395 251393 414429 251409
rect 414553 251469 414587 251485
rect 414553 251393 414587 251409
rect 414671 251469 414705 251485
rect 414671 251393 414705 251409
rect 414829 251469 414863 251485
rect 414829 251393 414863 251409
rect 414947 251469 414981 251485
rect 414947 251393 414981 251409
rect 415105 251469 415139 251485
rect 415105 251393 415139 251409
rect 415223 251469 415257 251485
rect 415223 251393 415257 251409
rect 415381 251469 415415 251485
rect 415381 251393 415415 251409
rect 415499 251469 415533 251485
rect 415499 251393 415533 251409
rect 415657 251469 415691 251485
rect 415657 251393 415691 251409
rect 415775 251469 415809 251485
rect 415775 251393 415809 251409
rect 415933 251469 415967 251485
rect 415933 251393 415967 251409
rect 416051 251469 416085 251485
rect 416051 251393 416085 251409
rect 416209 251469 416243 251485
rect 416209 251393 416243 251409
rect 416327 251469 416361 251485
rect 416327 251393 416361 251409
rect 416485 251469 416519 251485
rect 416485 251393 416519 251409
rect 416603 251469 416637 251485
rect 416603 251393 416637 251409
rect 416761 251469 416795 251485
rect 416761 251393 416795 251409
rect 416879 251469 416913 251485
rect 416879 251393 416913 251409
rect 417037 251469 417071 251485
rect 417037 251393 417071 251409
rect 417155 251469 417189 251485
rect 417155 251393 417189 251409
rect 417313 251469 417347 251485
rect 417313 251393 417347 251409
rect 417431 251469 417465 251485
rect 417431 251393 417465 251409
rect 417589 251469 417623 251485
rect 417589 251393 417623 251409
rect 417707 251469 417741 251485
rect 417707 251393 417741 251409
rect 417865 251469 417899 251485
rect 417865 251393 417899 251409
rect 417983 251469 418017 251485
rect 417983 251393 418017 251409
rect 418141 251469 418175 251485
rect 418141 251393 418175 251409
rect 418259 251469 418293 251485
rect 418259 251393 418293 251409
rect 418417 251469 418451 251485
rect 418417 251393 418451 251409
rect 418535 251469 418569 251485
rect 418535 251393 418569 251409
rect 418693 251469 418727 251485
rect 418693 251393 418727 251409
rect 418811 251469 418845 251485
rect 418811 251393 418845 251409
rect 418969 251469 419003 251485
rect 418969 251393 419003 251409
rect 419087 251469 419121 251485
rect 419087 251393 419121 251409
rect 419245 251469 419279 251485
rect 419245 251393 419279 251409
rect 419363 251469 419397 251485
rect 419363 251393 419397 251409
rect 419521 251469 419555 251485
rect 419521 251393 419555 251409
rect 419639 251469 419673 251485
rect 419639 251393 419673 251409
rect 419797 251469 419831 251485
rect 419797 251393 419831 251409
rect 419915 251469 419949 251485
rect 419915 251393 419949 251409
rect 420073 251469 420107 251485
rect 420073 251393 420107 251409
rect 420191 251469 420225 251485
rect 420191 251393 420225 251409
rect 420349 251469 420383 251485
rect 420349 251393 420383 251409
rect 420467 251469 420501 251485
rect 420467 251393 420501 251409
rect 420625 251469 420659 251485
rect 420625 251393 420659 251409
rect 420743 251469 420777 251485
rect 420743 251393 420777 251409
rect 420901 251469 420935 251485
rect 420901 251393 420935 251409
rect 421019 251469 421053 251485
rect 421019 251393 421053 251409
rect 421177 251469 421211 251485
rect 421177 251393 421211 251409
rect 421295 251469 421329 251485
rect 421295 251393 421329 251409
rect 421453 251469 421487 251485
rect 421453 251393 421487 251409
rect 421571 251469 421605 251485
rect 421571 251393 421605 251409
rect 421729 251469 421763 251485
rect 421729 251393 421763 251409
rect 421847 251469 421881 251485
rect 421847 251393 421881 251409
rect 422005 251469 422039 251485
rect 422005 251393 422039 251409
rect 422123 251469 422157 251485
rect 422123 251393 422157 251409
rect 422281 251469 422315 251485
rect 422281 251393 422315 251409
rect 422399 251469 422433 251485
rect 422399 251393 422433 251409
rect 422557 251469 422591 251485
rect 422557 251393 422591 251409
rect 422675 251469 422709 251485
rect 422675 251393 422709 251409
rect 422833 251469 422867 251485
rect 422833 251393 422867 251409
rect 422951 251469 422985 251485
rect 422951 251393 422985 251409
rect 423109 251469 423143 251485
rect 423109 251393 423143 251409
rect 423227 251469 423261 251485
rect 423227 251393 423261 251409
rect 423385 251469 423419 251485
rect 423385 251393 423419 251409
rect 423503 251469 423537 251485
rect 423503 251393 423537 251409
rect 423661 251469 423695 251485
rect 423661 251393 423695 251409
rect 423779 251469 423813 251485
rect 423779 251393 423813 251409
rect 423937 251469 423971 251485
rect 423937 251393 423971 251409
rect 424055 251469 424089 251485
rect 424055 251393 424089 251409
rect 424213 251469 424247 251485
rect 424213 251393 424247 251409
rect 424331 251469 424365 251485
rect 424331 251393 424365 251409
rect 424489 251469 424523 251485
rect 424489 251393 424523 251409
rect 424607 251469 424641 251485
rect 424607 251393 424641 251409
rect 424765 251469 424799 251485
rect 424765 251393 424799 251409
rect 424883 251469 424917 251485
rect 424883 251393 424917 251409
rect 425041 251469 425075 251485
rect 425041 251393 425075 251409
rect 425159 251469 425193 251485
rect 425159 251393 425193 251409
rect 425317 251469 425351 251485
rect 425317 251393 425351 251409
rect 425435 251469 425469 251485
rect 425435 251393 425469 251409
rect 425593 251469 425627 251485
rect 425593 251393 425627 251409
rect 425711 251469 425745 251485
rect 425711 251393 425745 251409
rect 425869 251469 425903 251485
rect 425869 251393 425903 251409
rect 425987 251469 426021 251485
rect 425987 251393 426021 251409
rect 426145 251469 426179 251485
rect 426145 251393 426179 251409
rect 426263 251469 426297 251485
rect 426263 251393 426297 251409
rect 426421 251469 426455 251485
rect 426421 251393 426455 251409
rect 426539 251469 426573 251485
rect 426539 251393 426573 251409
rect 426697 251469 426731 251485
rect 426697 251393 426731 251409
rect 426815 251469 426849 251485
rect 426815 251393 426849 251409
rect 426973 251469 427007 251485
rect 426973 251393 427007 251409
rect 427091 251469 427125 251485
rect 427091 251393 427125 251409
rect 427249 251469 427283 251485
rect 427249 251393 427283 251409
rect 234532 251314 238264 251370
rect 238342 251314 248751 251370
rect 413337 251325 413353 251359
rect 413421 251356 413437 251359
rect 413421 251325 413445 251356
rect 413613 251325 413629 251359
rect 413697 251325 413713 251359
rect 413889 251355 413905 251359
rect 413886 251325 413905 251355
rect 413973 251325 413989 251359
rect 414165 251351 414181 251359
rect 414162 251325 414181 251351
rect 414249 251325 414265 251359
rect 414441 251345 414457 251359
rect 414440 251325 414457 251345
rect 414525 251325 414541 251359
rect 414717 251341 414733 251359
rect 414716 251325 414733 251341
rect 414801 251325 414817 251359
rect 414993 251343 415009 251359
rect 414990 251325 415009 251343
rect 415077 251325 415093 251359
rect 415269 251341 415285 251359
rect 415268 251325 415285 251341
rect 415353 251325 415369 251359
rect 415545 251325 415561 251359
rect 415629 251325 415645 251359
rect 415821 251341 415837 251359
rect 415820 251325 415837 251341
rect 415905 251325 415921 251359
rect 416097 251325 416113 251359
rect 416181 251325 416197 251359
rect 416373 251351 416389 251359
rect 416370 251335 416389 251351
rect 416369 251325 416389 251335
rect 416457 251325 416473 251359
rect 416649 251351 416665 251359
rect 416646 251325 416665 251351
rect 416733 251325 416749 251359
rect 416925 251325 416941 251359
rect 417009 251325 417025 251359
rect 417201 251345 417217 251359
rect 417194 251325 417217 251345
rect 417285 251325 417301 251359
rect 417477 251325 417493 251359
rect 417561 251325 417577 251359
rect 417753 251345 417769 251359
rect 417752 251325 417769 251345
rect 417837 251325 417853 251359
rect 418029 251341 418045 251359
rect 418028 251325 418045 251341
rect 418113 251325 418129 251359
rect 418305 251349 418321 251359
rect 418302 251325 418321 251349
rect 418389 251325 418405 251359
rect 418581 251341 418597 251359
rect 418580 251325 418597 251341
rect 418665 251325 418681 251359
rect 418857 251343 418873 251359
rect 418850 251325 418873 251343
rect 418941 251325 418957 251359
rect 419133 251349 419149 251359
rect 419126 251325 419149 251349
rect 419217 251325 419233 251359
rect 419409 251355 419425 251359
rect 419408 251325 419425 251355
rect 419493 251325 419509 251359
rect 419685 251351 419701 251359
rect 419684 251325 419701 251351
rect 419769 251325 419785 251359
rect 419961 251351 419977 251359
rect 419958 251325 419977 251351
rect 420045 251325 420061 251359
rect 420237 251351 420253 251359
rect 420230 251325 420253 251351
rect 420321 251325 420337 251359
rect 420513 251351 420529 251359
rect 420512 251325 420529 251351
rect 420597 251325 420613 251359
rect 420789 251325 420805 251359
rect 420873 251325 420889 251359
rect 421065 251345 421081 251359
rect 421064 251325 421081 251345
rect 421149 251325 421165 251359
rect 421341 251325 421357 251359
rect 421425 251325 421441 251359
rect 421617 251325 421633 251359
rect 421701 251325 421717 251359
rect 421893 251337 421909 251359
rect 421886 251325 421909 251337
rect 421977 251325 421993 251359
rect 422169 251333 422185 251359
rect 422168 251325 422185 251333
rect 422253 251325 422269 251359
rect 422445 251325 422461 251359
rect 422529 251325 422545 251359
rect 422721 251333 422737 251359
rect 422720 251325 422737 251333
rect 422805 251325 422821 251359
rect 422997 251333 423013 251359
rect 422996 251325 423013 251333
rect 423081 251325 423097 251359
rect 423273 251349 423289 251359
rect 423266 251325 423289 251349
rect 423357 251325 423373 251359
rect 423549 251341 423565 251359
rect 423544 251325 423565 251341
rect 423633 251325 423649 251359
rect 423825 251325 423841 251359
rect 423909 251325 423925 251359
rect 424101 251325 424117 251359
rect 424185 251341 424201 251359
rect 424377 251345 424393 251359
rect 424185 251325 424206 251341
rect 234532 251303 248751 251314
rect 60236 251229 60270 251245
rect 59719 251208 60073 251210
rect 148668 251130 148784 251268
rect 234266 251252 234282 251294
rect 234336 251252 234346 251294
rect 234266 251232 234346 251252
rect 322693 251184 337190 251242
rect 148668 251086 148690 251130
rect 148762 251086 148784 251130
rect 148668 251060 148784 251086
rect 148726 251054 148784 251060
rect 322692 251144 337190 251184
rect 322692 250957 322779 251144
rect 322977 250957 323075 251144
rect 323253 250957 323351 251144
rect 323527 250957 323625 251144
rect 323805 250957 323903 251144
rect 324077 250957 324175 251144
rect 324355 250957 324453 251144
rect 324633 250957 324731 251144
rect 324911 250957 325009 251144
rect 325185 250957 325283 251144
rect 325461 250957 325559 251144
rect 325746 250957 325841 251144
rect 326015 250957 326113 251144
rect 326291 250957 326389 251144
rect 326563 250957 326661 251144
rect 326841 250957 326939 251144
rect 327113 250957 327211 251144
rect 327391 250957 327489 251144
rect 327667 250957 327765 251144
rect 322692 250934 322710 250957
rect 322694 250923 322710 250934
rect 322778 250923 322794 250957
rect 322970 250923 322986 250957
rect 323054 250933 323075 250957
rect 323054 250923 323070 250933
rect 323246 250923 323262 250957
rect 323330 250935 323351 250957
rect 323330 250923 323346 250935
rect 323522 250923 323538 250957
rect 323606 250931 323625 250957
rect 323606 250923 323622 250931
rect 323798 250923 323814 250957
rect 323882 250931 323903 250957
rect 323882 250923 323898 250931
rect 324074 250923 324090 250957
rect 324158 250933 324175 250957
rect 324158 250923 324174 250933
rect 324350 250923 324366 250957
rect 324434 250931 324453 250957
rect 324434 250923 324450 250931
rect 324626 250923 324642 250957
rect 324710 250931 324731 250957
rect 324710 250923 324726 250931
rect 324902 250923 324918 250957
rect 324986 250935 325009 250957
rect 324986 250923 325002 250935
rect 325178 250923 325194 250957
rect 325262 250931 325283 250957
rect 325262 250923 325278 250931
rect 325454 250923 325470 250957
rect 325538 250935 325559 250957
rect 325538 250923 325554 250935
rect 325730 250923 325746 250957
rect 325814 250934 325841 250957
rect 325814 250923 325830 250934
rect 326006 250923 326022 250957
rect 326090 250937 326113 250957
rect 326090 250923 326106 250937
rect 326282 250923 326298 250957
rect 326366 250927 326389 250957
rect 326366 250923 326382 250927
rect 326558 250923 326574 250957
rect 326642 250931 326661 250957
rect 326642 250923 326658 250931
rect 326834 250923 326850 250957
rect 326918 250931 326939 250957
rect 326918 250923 326934 250931
rect 327110 250923 327126 250957
rect 327194 250923 327211 250957
rect 327386 250923 327402 250957
rect 327470 250931 327489 250957
rect 327470 250923 327486 250931
rect 327662 250923 327678 250957
rect 327746 250931 327765 250957
rect 327937 250957 328035 251144
rect 328223 250957 328321 251144
rect 328495 250957 328593 251144
rect 328775 250957 328873 251144
rect 329049 250957 329147 251144
rect 329601 250957 329699 251144
rect 329877 250957 329975 251144
rect 330153 250957 330251 251144
rect 330429 250957 330527 251144
rect 330705 250957 330803 251144
rect 330981 250957 331079 251144
rect 331259 250957 331357 251144
rect 331535 250957 331633 251144
rect 331807 250957 331905 251144
rect 332085 250957 332183 251144
rect 332361 250957 332459 251144
rect 332639 250957 332737 251144
rect 332913 250957 333011 251144
rect 333189 250957 333287 251144
rect 333467 250957 333565 251144
rect 333743 250957 333841 251144
rect 334019 250957 334117 251144
rect 334295 250957 334393 251144
rect 334571 250957 334669 251144
rect 334845 250957 334943 251144
rect 335125 250957 335223 251144
rect 335401 250957 335499 251144
rect 335673 250957 335771 251144
rect 335949 250957 336047 251144
rect 336219 250957 336317 251144
rect 336511 250957 336609 251144
rect 327746 250923 327762 250931
rect 327937 250929 327954 250957
rect 327938 250923 327954 250929
rect 328022 250923 328038 250957
rect 328214 250923 328230 250957
rect 328298 250927 328321 250957
rect 328298 250923 328314 250927
rect 328490 250923 328506 250957
rect 328574 250927 328593 250957
rect 328574 250923 328590 250927
rect 328766 250923 328782 250957
rect 328850 250927 328873 250957
rect 328850 250923 328866 250927
rect 329042 250923 329058 250957
rect 329126 250927 329147 250957
rect 329126 250923 329142 250927
rect 329318 250923 329334 250957
rect 329402 250923 329418 250957
rect 329594 250923 329610 250957
rect 329678 250927 329699 250957
rect 329678 250923 329694 250927
rect 329870 250923 329886 250957
rect 329954 250929 329975 250957
rect 329954 250923 329970 250929
rect 330146 250923 330162 250957
rect 330230 250929 330251 250957
rect 330230 250923 330246 250929
rect 330422 250923 330438 250957
rect 330506 250931 330527 250957
rect 330506 250923 330522 250931
rect 330698 250923 330714 250957
rect 330782 250929 330803 250957
rect 330782 250923 330798 250929
rect 330974 250923 330990 250957
rect 331058 250929 331079 250957
rect 331058 250923 331074 250929
rect 331250 250923 331266 250957
rect 331334 250929 331357 250957
rect 331334 250923 331350 250929
rect 331526 250923 331542 250957
rect 331610 250929 331633 250957
rect 331610 250923 331626 250929
rect 331802 250923 331818 250957
rect 331886 250927 331905 250957
rect 331886 250923 331902 250927
rect 332078 250923 332094 250957
rect 332162 250927 332183 250957
rect 332162 250923 332178 250927
rect 332354 250923 332370 250957
rect 332438 250931 332459 250957
rect 332438 250923 332454 250931
rect 332630 250923 332646 250957
rect 332714 250933 332737 250957
rect 332714 250923 332730 250933
rect 332906 250923 332922 250957
rect 332990 250929 333011 250957
rect 332990 250923 333006 250929
rect 333182 250923 333198 250957
rect 333266 250933 333287 250957
rect 333266 250923 333282 250933
rect 333458 250923 333474 250957
rect 333542 250933 333565 250957
rect 333542 250923 333558 250933
rect 333734 250923 333750 250957
rect 333818 250935 333841 250957
rect 333818 250923 333834 250935
rect 334010 250923 334026 250957
rect 334094 250931 334117 250957
rect 334094 250923 334110 250931
rect 334286 250923 334302 250957
rect 334370 250933 334393 250957
rect 334370 250923 334386 250933
rect 334562 250923 334578 250957
rect 334646 250933 334669 250957
rect 334646 250923 334662 250933
rect 334838 250923 334854 250957
rect 334922 250935 334943 250957
rect 334922 250923 334938 250935
rect 335114 250923 335130 250957
rect 335198 250935 335223 250957
rect 335198 250923 335214 250935
rect 335390 250923 335406 250957
rect 335474 250935 335499 250957
rect 335474 250923 335490 250935
rect 335666 250923 335682 250957
rect 335750 250935 335771 250957
rect 335750 250923 335766 250935
rect 335942 250923 335958 250957
rect 336026 250925 336047 250957
rect 336026 250923 336042 250925
rect 336218 250923 336234 250957
rect 336302 250923 336318 250957
rect 336494 250923 336510 250957
rect 336578 250925 336609 250957
rect 336740 250999 336774 251015
rect 336578 250923 336594 250925
rect 322648 250873 322682 250889
rect 322648 250797 322682 250813
rect 322806 250873 322840 250889
rect 322806 250797 322840 250813
rect 322924 250873 322958 250889
rect 322924 250797 322958 250813
rect 323082 250873 323116 250889
rect 323082 250797 323116 250813
rect 323200 250873 323234 250889
rect 323200 250797 323234 250813
rect 323358 250873 323392 250889
rect 323358 250797 323392 250813
rect 323476 250873 323510 250889
rect 323476 250797 323510 250813
rect 323634 250873 323668 250889
rect 323634 250797 323668 250813
rect 323752 250873 323786 250889
rect 323752 250797 323786 250813
rect 323910 250873 323944 250889
rect 323910 250797 323944 250813
rect 324028 250873 324062 250889
rect 324028 250797 324062 250813
rect 324186 250873 324220 250889
rect 324186 250797 324220 250813
rect 324304 250873 324338 250889
rect 324304 250797 324338 250813
rect 324462 250873 324496 250889
rect 324462 250797 324496 250813
rect 324580 250873 324614 250889
rect 324580 250797 324614 250813
rect 324738 250873 324772 250889
rect 324738 250797 324772 250813
rect 324856 250873 324890 250889
rect 324856 250797 324890 250813
rect 325014 250873 325048 250889
rect 325014 250797 325048 250813
rect 325132 250873 325166 250889
rect 325132 250797 325166 250813
rect 325290 250873 325324 250889
rect 325290 250797 325324 250813
rect 325408 250873 325442 250889
rect 325408 250797 325442 250813
rect 325566 250873 325600 250889
rect 325566 250797 325600 250813
rect 325684 250873 325718 250889
rect 325684 250797 325718 250813
rect 325842 250873 325876 250889
rect 325842 250797 325876 250813
rect 325960 250873 325994 250889
rect 325960 250797 325994 250813
rect 326118 250873 326152 250889
rect 326118 250797 326152 250813
rect 326236 250873 326270 250889
rect 326236 250797 326270 250813
rect 326394 250873 326428 250889
rect 326394 250797 326428 250813
rect 326512 250873 326546 250889
rect 326512 250797 326546 250813
rect 326670 250873 326704 250889
rect 326670 250797 326704 250813
rect 326788 250873 326822 250889
rect 326788 250797 326822 250813
rect 326946 250873 326980 250889
rect 326946 250797 326980 250813
rect 327064 250873 327098 250889
rect 327064 250797 327098 250813
rect 327222 250873 327256 250889
rect 327222 250797 327256 250813
rect 327340 250873 327374 250889
rect 327340 250797 327374 250813
rect 327498 250873 327532 250889
rect 327498 250797 327532 250813
rect 327616 250873 327650 250889
rect 327616 250797 327650 250813
rect 327774 250873 327808 250889
rect 327774 250797 327808 250813
rect 327892 250873 327926 250889
rect 327892 250797 327926 250813
rect 328050 250873 328084 250889
rect 328050 250797 328084 250813
rect 328168 250873 328202 250889
rect 328168 250797 328202 250813
rect 328326 250873 328360 250889
rect 328326 250797 328360 250813
rect 328444 250873 328478 250889
rect 328444 250797 328478 250813
rect 328602 250873 328636 250889
rect 328602 250797 328636 250813
rect 328720 250873 328754 250889
rect 328720 250797 328754 250813
rect 328878 250873 328912 250889
rect 328878 250797 328912 250813
rect 328996 250873 329030 250889
rect 328996 250797 329030 250813
rect 329154 250873 329188 250889
rect 329154 250797 329188 250813
rect 329272 250873 329306 250889
rect 329272 250797 329306 250813
rect 329430 250873 329464 250889
rect 329430 250797 329464 250813
rect 329548 250873 329582 250889
rect 329548 250797 329582 250813
rect 329706 250873 329740 250889
rect 329706 250797 329740 250813
rect 329824 250873 329858 250889
rect 329824 250797 329858 250813
rect 329982 250873 330016 250889
rect 329982 250797 330016 250813
rect 330100 250873 330134 250889
rect 330100 250797 330134 250813
rect 330258 250873 330292 250889
rect 330258 250797 330292 250813
rect 330376 250873 330410 250889
rect 330376 250797 330410 250813
rect 330534 250873 330568 250889
rect 330534 250797 330568 250813
rect 330652 250873 330686 250889
rect 330652 250797 330686 250813
rect 330810 250873 330844 250889
rect 330810 250797 330844 250813
rect 330928 250873 330962 250889
rect 330928 250797 330962 250813
rect 331086 250873 331120 250889
rect 331086 250797 331120 250813
rect 331204 250873 331238 250889
rect 331204 250797 331238 250813
rect 331362 250873 331396 250889
rect 331362 250797 331396 250813
rect 331480 250873 331514 250889
rect 331480 250797 331514 250813
rect 331638 250873 331672 250889
rect 331638 250797 331672 250813
rect 331756 250873 331790 250889
rect 331756 250797 331790 250813
rect 331914 250873 331948 250889
rect 331914 250797 331948 250813
rect 332032 250873 332066 250889
rect 332032 250797 332066 250813
rect 332190 250873 332224 250889
rect 332190 250797 332224 250813
rect 332308 250873 332342 250889
rect 332308 250797 332342 250813
rect 332466 250873 332500 250889
rect 332466 250797 332500 250813
rect 332584 250873 332618 250889
rect 332584 250797 332618 250813
rect 332742 250873 332776 250889
rect 332742 250797 332776 250813
rect 332860 250873 332894 250889
rect 332860 250797 332894 250813
rect 333018 250873 333052 250889
rect 333018 250797 333052 250813
rect 333136 250873 333170 250889
rect 333136 250797 333170 250813
rect 333294 250873 333328 250889
rect 333294 250797 333328 250813
rect 333412 250873 333446 250889
rect 333412 250797 333446 250813
rect 333570 250873 333604 250889
rect 333570 250797 333604 250813
rect 333688 250873 333722 250889
rect 333688 250797 333722 250813
rect 333846 250873 333880 250889
rect 333846 250797 333880 250813
rect 333964 250873 333998 250889
rect 333964 250797 333998 250813
rect 334122 250873 334156 250889
rect 334122 250797 334156 250813
rect 334240 250873 334274 250889
rect 334240 250797 334274 250813
rect 334398 250873 334432 250889
rect 334398 250797 334432 250813
rect 334516 250873 334550 250889
rect 334516 250797 334550 250813
rect 334674 250873 334708 250889
rect 334674 250797 334708 250813
rect 334792 250873 334826 250889
rect 334792 250797 334826 250813
rect 334950 250873 334984 250889
rect 334950 250797 334984 250813
rect 335068 250873 335102 250889
rect 335068 250797 335102 250813
rect 335226 250873 335260 250889
rect 335226 250797 335260 250813
rect 335344 250873 335378 250889
rect 335344 250797 335378 250813
rect 335502 250873 335536 250889
rect 335502 250797 335536 250813
rect 335620 250873 335654 250889
rect 335620 250797 335654 250813
rect 335778 250873 335812 250889
rect 335778 250797 335812 250813
rect 335896 250873 335930 250889
rect 335896 250797 335930 250813
rect 336054 250873 336088 250889
rect 336054 250797 336088 250813
rect 336172 250873 336206 250889
rect 336172 250797 336206 250813
rect 336330 250873 336364 250889
rect 336330 250797 336364 250813
rect 336448 250873 336482 250889
rect 336448 250797 336482 250813
rect 336606 250873 336640 250889
rect 336606 250797 336640 250813
rect 322694 250729 322710 250763
rect 322778 250760 322794 250763
rect 322778 250729 322802 250760
rect 322970 250729 322986 250763
rect 323054 250729 323070 250763
rect 323246 250759 323262 250763
rect 323243 250729 323262 250759
rect 323330 250729 323346 250763
rect 323522 250755 323538 250763
rect 323519 250729 323538 250755
rect 323606 250729 323622 250763
rect 323798 250749 323814 250763
rect 323797 250729 323814 250749
rect 323882 250729 323898 250763
rect 324074 250745 324090 250763
rect 324073 250729 324090 250745
rect 324158 250729 324174 250763
rect 324350 250747 324366 250763
rect 324347 250729 324366 250747
rect 324434 250729 324450 250763
rect 324626 250745 324642 250763
rect 324625 250729 324642 250745
rect 324710 250729 324726 250763
rect 324902 250729 324918 250763
rect 324986 250729 325002 250763
rect 325178 250745 325194 250763
rect 325177 250729 325194 250745
rect 325262 250729 325278 250763
rect 325454 250729 325470 250763
rect 325538 250729 325554 250763
rect 325730 250755 325746 250763
rect 325727 250739 325746 250755
rect 325726 250729 325746 250739
rect 325814 250729 325830 250763
rect 326006 250755 326022 250763
rect 326003 250729 326022 250755
rect 326090 250729 326106 250763
rect 326282 250729 326298 250763
rect 326366 250729 326382 250763
rect 326558 250749 326574 250763
rect 326551 250729 326574 250749
rect 326642 250729 326658 250763
rect 326834 250729 326850 250763
rect 326918 250729 326934 250763
rect 327110 250749 327126 250763
rect 327109 250729 327126 250749
rect 327194 250729 327210 250763
rect 327386 250745 327402 250763
rect 327385 250729 327402 250745
rect 327470 250729 327486 250763
rect 327662 250753 327678 250763
rect 327659 250729 327678 250753
rect 327746 250729 327762 250763
rect 327938 250745 327954 250763
rect 327937 250729 327954 250745
rect 328022 250729 328038 250763
rect 328214 250747 328230 250763
rect 328207 250729 328230 250747
rect 328298 250729 328314 250763
rect 328490 250753 328506 250763
rect 328483 250729 328506 250753
rect 328574 250729 328590 250763
rect 328766 250759 328782 250763
rect 328765 250729 328782 250759
rect 328850 250729 328866 250763
rect 329042 250755 329058 250763
rect 329041 250729 329058 250755
rect 329126 250729 329142 250763
rect 329318 250755 329334 250763
rect 329315 250729 329334 250755
rect 329402 250729 329418 250763
rect 329594 250755 329610 250763
rect 329587 250729 329610 250755
rect 329678 250729 329694 250763
rect 329870 250755 329886 250763
rect 329869 250729 329886 250755
rect 329954 250729 329970 250763
rect 330146 250729 330162 250763
rect 330230 250729 330246 250763
rect 330422 250749 330438 250763
rect 330421 250729 330438 250749
rect 330506 250729 330522 250763
rect 330698 250729 330714 250763
rect 330782 250729 330798 250763
rect 330974 250729 330990 250763
rect 331058 250729 331074 250763
rect 331250 250741 331266 250763
rect 331243 250729 331266 250741
rect 331334 250729 331350 250763
rect 331526 250737 331542 250763
rect 331525 250729 331542 250737
rect 331610 250729 331626 250763
rect 331802 250729 331818 250763
rect 331886 250729 331902 250763
rect 332078 250737 332094 250763
rect 332077 250729 332094 250737
rect 332162 250729 332178 250763
rect 332354 250737 332370 250763
rect 332353 250729 332370 250737
rect 332438 250729 332454 250763
rect 332630 250753 332646 250763
rect 332623 250729 332646 250753
rect 332714 250729 332730 250763
rect 332906 250745 332922 250763
rect 332901 250729 332922 250745
rect 332990 250729 333006 250763
rect 333182 250729 333198 250763
rect 333266 250729 333282 250763
rect 333458 250729 333474 250763
rect 333542 250745 333558 250763
rect 333734 250749 333750 250763
rect 333542 250729 333563 250745
rect 322700 250520 322802 250729
rect 322971 250520 323069 250729
rect 323243 250520 323341 250729
rect 323519 250520 323617 250729
rect 323797 250520 323895 250729
rect 324073 250520 324171 250729
rect 324347 250520 324445 250729
rect 324625 250520 324723 250729
rect 324903 250520 325001 250729
rect 325177 250520 325275 250729
rect 325455 250520 325553 250729
rect 325726 250520 325826 250729
rect 326003 250520 326101 250729
rect 326283 250520 326381 250729
rect 326551 250520 326649 250729
rect 326835 250520 326933 250729
rect 327109 250520 327207 250729
rect 327385 250520 327483 250729
rect 327659 250520 327757 250729
rect 327937 250520 328035 250729
rect 328207 250520 328305 250729
rect 328483 250520 328581 250729
rect 328765 250520 328863 250729
rect 329041 250520 329139 250729
rect 329315 250714 329413 250729
rect 329587 250520 329685 250729
rect 329869 250520 329967 250729
rect 330147 250520 330245 250729
rect 330421 250520 330519 250729
rect 330699 250520 330797 250729
rect 330975 250520 331073 250729
rect 331243 250520 331341 250729
rect 331525 250520 331623 250729
rect 331803 250520 331901 250729
rect 332077 250520 332175 250729
rect 332353 250520 332451 250729
rect 332623 250520 332721 250729
rect 332901 250520 332999 250729
rect 333183 250520 333281 250729
rect 333465 250520 333563 250729
rect 333733 250729 333750 250749
rect 333818 250729 333834 250763
rect 334010 250749 334026 250763
rect 334009 250729 334026 250749
rect 334094 250729 334110 250763
rect 334286 250749 334302 250763
rect 334279 250729 334302 250749
rect 334370 250729 334386 250763
rect 334562 250755 334578 250763
rect 334557 250729 334578 250755
rect 334646 250729 334662 250763
rect 334838 250729 334854 250763
rect 334922 250729 334938 250763
rect 335114 250729 335130 250763
rect 335198 250755 335214 250763
rect 335198 250729 335217 250755
rect 335390 250753 335406 250763
rect 333733 250520 333831 250729
rect 334009 250520 334107 250729
rect 334279 250520 334377 250729
rect 334557 250520 334655 250729
rect 334839 250520 334937 250729
rect 335119 250520 335217 250729
rect 335385 250729 335406 250753
rect 335474 250729 335490 250763
rect 335666 250747 335682 250763
rect 335661 250729 335682 250747
rect 335750 250729 335766 250763
rect 335942 250753 335958 250763
rect 335941 250729 335958 250753
rect 336026 250729 336042 250763
rect 336218 250729 336234 250763
rect 336302 250753 336318 250763
rect 336302 250729 336323 250753
rect 336494 250729 336510 250763
rect 336578 250757 336594 250763
rect 336578 250729 336601 250757
rect 335385 250520 335483 250729
rect 335661 250520 335759 250729
rect 335941 250520 336039 250729
rect 336225 250520 336323 250729
rect 336503 250520 336601 250729
rect 336740 250671 336774 250687
rect 337092 250520 337190 251144
rect 413343 251116 413445 251325
rect 413614 251116 413712 251325
rect 413886 251116 413984 251325
rect 414162 251116 414260 251325
rect 414440 251116 414538 251325
rect 414716 251116 414814 251325
rect 414990 251116 415088 251325
rect 415268 251116 415366 251325
rect 415546 251116 415644 251325
rect 415820 251116 415918 251325
rect 416098 251116 416196 251325
rect 416369 251116 416469 251325
rect 416646 251116 416744 251325
rect 416926 251116 417024 251325
rect 417194 251116 417292 251325
rect 417478 251116 417576 251325
rect 417752 251116 417850 251325
rect 418028 251116 418126 251325
rect 418302 251116 418400 251325
rect 418580 251116 418678 251325
rect 418850 251116 418948 251325
rect 419126 251116 419224 251325
rect 419408 251116 419506 251325
rect 419684 251116 419782 251325
rect 419958 251310 420056 251325
rect 420230 251116 420328 251325
rect 420512 251116 420610 251325
rect 420790 251116 420888 251325
rect 421064 251116 421162 251325
rect 421342 251116 421440 251325
rect 421618 251116 421716 251325
rect 421886 251116 421984 251325
rect 422168 251116 422266 251325
rect 422446 251116 422544 251325
rect 422720 251116 422818 251325
rect 422996 251116 423094 251325
rect 423266 251116 423364 251325
rect 423544 251116 423642 251325
rect 423826 251116 423924 251325
rect 424108 251116 424206 251325
rect 424376 251325 424393 251345
rect 424461 251325 424477 251359
rect 424653 251345 424669 251359
rect 424652 251325 424669 251345
rect 424737 251325 424753 251359
rect 424929 251345 424945 251359
rect 424922 251325 424945 251345
rect 425013 251325 425029 251359
rect 425205 251351 425221 251359
rect 425200 251325 425221 251351
rect 425289 251325 425305 251359
rect 425481 251325 425497 251359
rect 425565 251325 425581 251359
rect 425757 251325 425773 251359
rect 425841 251351 425857 251359
rect 425841 251325 425860 251351
rect 426033 251349 426049 251359
rect 424376 251116 424474 251325
rect 424652 251116 424750 251325
rect 424922 251116 425020 251325
rect 425200 251116 425298 251325
rect 425482 251116 425580 251325
rect 425762 251116 425860 251325
rect 426028 251325 426049 251349
rect 426117 251325 426133 251359
rect 426309 251343 426325 251359
rect 426304 251325 426325 251343
rect 426393 251325 426409 251359
rect 426585 251349 426601 251359
rect 426584 251325 426601 251349
rect 426669 251325 426685 251359
rect 426861 251325 426877 251359
rect 426945 251349 426961 251359
rect 426945 251325 426966 251349
rect 427137 251325 427153 251359
rect 427221 251353 427237 251359
rect 427221 251325 427244 251353
rect 426028 251116 426126 251325
rect 426304 251116 426402 251325
rect 426584 251116 426682 251325
rect 426868 251116 426966 251325
rect 427146 251116 427244 251325
rect 427383 251267 427417 251283
rect 427735 251116 427833 251740
rect 503335 251740 517833 251780
rect 503335 251553 503422 251740
rect 503620 251553 503718 251740
rect 503896 251553 503994 251740
rect 504170 251553 504268 251740
rect 504448 251553 504546 251740
rect 504720 251553 504818 251740
rect 504998 251553 505096 251740
rect 505276 251553 505374 251740
rect 505554 251553 505652 251740
rect 505828 251553 505926 251740
rect 506104 251553 506202 251740
rect 506389 251553 506484 251740
rect 506658 251553 506756 251740
rect 506934 251553 507032 251740
rect 507206 251553 507304 251740
rect 507484 251553 507582 251740
rect 507756 251553 507854 251740
rect 508034 251553 508132 251740
rect 508310 251553 508408 251740
rect 503335 251530 503353 251553
rect 503337 251519 503353 251530
rect 503421 251519 503437 251553
rect 503613 251519 503629 251553
rect 503697 251529 503718 251553
rect 503697 251519 503713 251529
rect 503889 251519 503905 251553
rect 503973 251531 503994 251553
rect 503973 251519 503989 251531
rect 504165 251519 504181 251553
rect 504249 251527 504268 251553
rect 504249 251519 504265 251527
rect 504441 251519 504457 251553
rect 504525 251527 504546 251553
rect 504525 251519 504541 251527
rect 504717 251519 504733 251553
rect 504801 251529 504818 251553
rect 504801 251519 504817 251529
rect 504993 251519 505009 251553
rect 505077 251527 505096 251553
rect 505077 251519 505093 251527
rect 505269 251519 505285 251553
rect 505353 251527 505374 251553
rect 505353 251519 505369 251527
rect 505545 251519 505561 251553
rect 505629 251531 505652 251553
rect 505629 251519 505645 251531
rect 505821 251519 505837 251553
rect 505905 251527 505926 251553
rect 505905 251519 505921 251527
rect 506097 251519 506113 251553
rect 506181 251531 506202 251553
rect 506181 251519 506197 251531
rect 506373 251519 506389 251553
rect 506457 251530 506484 251553
rect 506457 251519 506473 251530
rect 506649 251519 506665 251553
rect 506733 251533 506756 251553
rect 506733 251519 506749 251533
rect 506925 251519 506941 251553
rect 507009 251523 507032 251553
rect 507009 251519 507025 251523
rect 507201 251519 507217 251553
rect 507285 251527 507304 251553
rect 507285 251519 507301 251527
rect 507477 251519 507493 251553
rect 507561 251527 507582 251553
rect 507561 251519 507577 251527
rect 507753 251519 507769 251553
rect 507837 251519 507854 251553
rect 508029 251519 508045 251553
rect 508113 251527 508132 251553
rect 508113 251519 508129 251527
rect 508305 251519 508321 251553
rect 508389 251527 508408 251553
rect 508580 251553 508678 251740
rect 508866 251553 508964 251740
rect 509138 251553 509236 251740
rect 509418 251553 509516 251740
rect 509692 251553 509790 251740
rect 510244 251553 510342 251740
rect 510520 251553 510618 251740
rect 510796 251553 510894 251740
rect 511072 251553 511170 251740
rect 511348 251553 511446 251740
rect 511624 251553 511722 251740
rect 511902 251553 512000 251740
rect 512178 251553 512276 251740
rect 512450 251553 512548 251740
rect 512728 251553 512826 251740
rect 513004 251553 513102 251740
rect 513282 251553 513380 251740
rect 513556 251553 513654 251740
rect 513832 251553 513930 251740
rect 514110 251553 514208 251740
rect 514386 251553 514484 251740
rect 514662 251553 514760 251740
rect 514938 251553 515036 251740
rect 515214 251553 515312 251740
rect 515488 251553 515586 251740
rect 515768 251553 515866 251740
rect 516044 251553 516142 251740
rect 516316 251553 516414 251740
rect 516592 251553 516690 251740
rect 516862 251553 516960 251740
rect 517154 251553 517252 251740
rect 508389 251519 508405 251527
rect 508580 251525 508597 251553
rect 508581 251519 508597 251525
rect 508665 251519 508681 251553
rect 508857 251519 508873 251553
rect 508941 251523 508964 251553
rect 508941 251519 508957 251523
rect 509133 251519 509149 251553
rect 509217 251523 509236 251553
rect 509217 251519 509233 251523
rect 509409 251519 509425 251553
rect 509493 251523 509516 251553
rect 509493 251519 509509 251523
rect 509685 251519 509701 251553
rect 509769 251523 509790 251553
rect 509769 251519 509785 251523
rect 509961 251519 509977 251553
rect 510045 251519 510061 251553
rect 510237 251519 510253 251553
rect 510321 251523 510342 251553
rect 510321 251519 510337 251523
rect 510513 251519 510529 251553
rect 510597 251525 510618 251553
rect 510597 251519 510613 251525
rect 510789 251519 510805 251553
rect 510873 251525 510894 251553
rect 510873 251519 510889 251525
rect 511065 251519 511081 251553
rect 511149 251527 511170 251553
rect 511149 251519 511165 251527
rect 511341 251519 511357 251553
rect 511425 251525 511446 251553
rect 511425 251519 511441 251525
rect 511617 251519 511633 251553
rect 511701 251525 511722 251553
rect 511701 251519 511717 251525
rect 511893 251519 511909 251553
rect 511977 251525 512000 251553
rect 511977 251519 511993 251525
rect 512169 251519 512185 251553
rect 512253 251525 512276 251553
rect 512253 251519 512269 251525
rect 512445 251519 512461 251553
rect 512529 251523 512548 251553
rect 512529 251519 512545 251523
rect 512721 251519 512737 251553
rect 512805 251523 512826 251553
rect 512805 251519 512821 251523
rect 512997 251519 513013 251553
rect 513081 251527 513102 251553
rect 513081 251519 513097 251527
rect 513273 251519 513289 251553
rect 513357 251529 513380 251553
rect 513357 251519 513373 251529
rect 513549 251519 513565 251553
rect 513633 251525 513654 251553
rect 513633 251519 513649 251525
rect 513825 251519 513841 251553
rect 513909 251529 513930 251553
rect 513909 251519 513925 251529
rect 514101 251519 514117 251553
rect 514185 251529 514208 251553
rect 514185 251519 514201 251529
rect 514377 251519 514393 251553
rect 514461 251531 514484 251553
rect 514461 251519 514477 251531
rect 514653 251519 514669 251553
rect 514737 251527 514760 251553
rect 514737 251519 514753 251527
rect 514929 251519 514945 251553
rect 515013 251529 515036 251553
rect 515013 251519 515029 251529
rect 515205 251519 515221 251553
rect 515289 251529 515312 251553
rect 515289 251519 515305 251529
rect 515481 251519 515497 251553
rect 515565 251531 515586 251553
rect 515565 251519 515581 251531
rect 515757 251519 515773 251553
rect 515841 251531 515866 251553
rect 515841 251519 515857 251531
rect 516033 251519 516049 251553
rect 516117 251531 516142 251553
rect 516117 251519 516133 251531
rect 516309 251519 516325 251553
rect 516393 251531 516414 251553
rect 516393 251519 516409 251531
rect 516585 251519 516601 251553
rect 516669 251521 516690 251553
rect 516669 251519 516685 251521
rect 516861 251519 516877 251553
rect 516945 251519 516961 251553
rect 517137 251519 517153 251553
rect 517221 251521 517252 251553
rect 517383 251595 517417 251611
rect 517221 251519 517237 251521
rect 503291 251469 503325 251485
rect 503291 251393 503325 251409
rect 503449 251469 503483 251485
rect 503449 251393 503483 251409
rect 503567 251469 503601 251485
rect 503567 251393 503601 251409
rect 503725 251469 503759 251485
rect 503725 251393 503759 251409
rect 503843 251469 503877 251485
rect 503843 251393 503877 251409
rect 504001 251469 504035 251485
rect 504001 251393 504035 251409
rect 504119 251469 504153 251485
rect 504119 251393 504153 251409
rect 504277 251469 504311 251485
rect 504277 251393 504311 251409
rect 504395 251469 504429 251485
rect 504395 251393 504429 251409
rect 504553 251469 504587 251485
rect 504553 251393 504587 251409
rect 504671 251469 504705 251485
rect 504671 251393 504705 251409
rect 504829 251469 504863 251485
rect 504829 251393 504863 251409
rect 504947 251469 504981 251485
rect 504947 251393 504981 251409
rect 505105 251469 505139 251485
rect 505105 251393 505139 251409
rect 505223 251469 505257 251485
rect 505223 251393 505257 251409
rect 505381 251469 505415 251485
rect 505381 251393 505415 251409
rect 505499 251469 505533 251485
rect 505499 251393 505533 251409
rect 505657 251469 505691 251485
rect 505657 251393 505691 251409
rect 505775 251469 505809 251485
rect 505775 251393 505809 251409
rect 505933 251469 505967 251485
rect 505933 251393 505967 251409
rect 506051 251469 506085 251485
rect 506051 251393 506085 251409
rect 506209 251469 506243 251485
rect 506209 251393 506243 251409
rect 506327 251469 506361 251485
rect 506327 251393 506361 251409
rect 506485 251469 506519 251485
rect 506485 251393 506519 251409
rect 506603 251469 506637 251485
rect 506603 251393 506637 251409
rect 506761 251469 506795 251485
rect 506761 251393 506795 251409
rect 506879 251469 506913 251485
rect 506879 251393 506913 251409
rect 507037 251469 507071 251485
rect 507037 251393 507071 251409
rect 507155 251469 507189 251485
rect 507155 251393 507189 251409
rect 507313 251469 507347 251485
rect 507313 251393 507347 251409
rect 507431 251469 507465 251485
rect 507431 251393 507465 251409
rect 507589 251469 507623 251485
rect 507589 251393 507623 251409
rect 507707 251469 507741 251485
rect 507707 251393 507741 251409
rect 507865 251469 507899 251485
rect 507865 251393 507899 251409
rect 507983 251469 508017 251485
rect 507983 251393 508017 251409
rect 508141 251469 508175 251485
rect 508141 251393 508175 251409
rect 508259 251469 508293 251485
rect 508259 251393 508293 251409
rect 508417 251469 508451 251485
rect 508417 251393 508451 251409
rect 508535 251469 508569 251485
rect 508535 251393 508569 251409
rect 508693 251469 508727 251485
rect 508693 251393 508727 251409
rect 508811 251469 508845 251485
rect 508811 251393 508845 251409
rect 508969 251469 509003 251485
rect 508969 251393 509003 251409
rect 509087 251469 509121 251485
rect 509087 251393 509121 251409
rect 509245 251469 509279 251485
rect 509245 251393 509279 251409
rect 509363 251469 509397 251485
rect 509363 251393 509397 251409
rect 509521 251469 509555 251485
rect 509521 251393 509555 251409
rect 509639 251469 509673 251485
rect 509639 251393 509673 251409
rect 509797 251469 509831 251485
rect 509797 251393 509831 251409
rect 509915 251469 509949 251485
rect 509915 251393 509949 251409
rect 510073 251469 510107 251485
rect 510073 251393 510107 251409
rect 510191 251469 510225 251485
rect 510191 251393 510225 251409
rect 510349 251469 510383 251485
rect 510349 251393 510383 251409
rect 510467 251469 510501 251485
rect 510467 251393 510501 251409
rect 510625 251469 510659 251485
rect 510625 251393 510659 251409
rect 510743 251469 510777 251485
rect 510743 251393 510777 251409
rect 510901 251469 510935 251485
rect 510901 251393 510935 251409
rect 511019 251469 511053 251485
rect 511019 251393 511053 251409
rect 511177 251469 511211 251485
rect 511177 251393 511211 251409
rect 511295 251469 511329 251485
rect 511295 251393 511329 251409
rect 511453 251469 511487 251485
rect 511453 251393 511487 251409
rect 511571 251469 511605 251485
rect 511571 251393 511605 251409
rect 511729 251469 511763 251485
rect 511729 251393 511763 251409
rect 511847 251469 511881 251485
rect 511847 251393 511881 251409
rect 512005 251469 512039 251485
rect 512005 251393 512039 251409
rect 512123 251469 512157 251485
rect 512123 251393 512157 251409
rect 512281 251469 512315 251485
rect 512281 251393 512315 251409
rect 512399 251469 512433 251485
rect 512399 251393 512433 251409
rect 512557 251469 512591 251485
rect 512557 251393 512591 251409
rect 512675 251469 512709 251485
rect 512675 251393 512709 251409
rect 512833 251469 512867 251485
rect 512833 251393 512867 251409
rect 512951 251469 512985 251485
rect 512951 251393 512985 251409
rect 513109 251469 513143 251485
rect 513109 251393 513143 251409
rect 513227 251469 513261 251485
rect 513227 251393 513261 251409
rect 513385 251469 513419 251485
rect 513385 251393 513419 251409
rect 513503 251469 513537 251485
rect 513503 251393 513537 251409
rect 513661 251469 513695 251485
rect 513661 251393 513695 251409
rect 513779 251469 513813 251485
rect 513779 251393 513813 251409
rect 513937 251469 513971 251485
rect 513937 251393 513971 251409
rect 514055 251469 514089 251485
rect 514055 251393 514089 251409
rect 514213 251469 514247 251485
rect 514213 251393 514247 251409
rect 514331 251469 514365 251485
rect 514331 251393 514365 251409
rect 514489 251469 514523 251485
rect 514489 251393 514523 251409
rect 514607 251469 514641 251485
rect 514607 251393 514641 251409
rect 514765 251469 514799 251485
rect 514765 251393 514799 251409
rect 514883 251469 514917 251485
rect 514883 251393 514917 251409
rect 515041 251469 515075 251485
rect 515041 251393 515075 251409
rect 515159 251469 515193 251485
rect 515159 251393 515193 251409
rect 515317 251469 515351 251485
rect 515317 251393 515351 251409
rect 515435 251469 515469 251485
rect 515435 251393 515469 251409
rect 515593 251469 515627 251485
rect 515593 251393 515627 251409
rect 515711 251469 515745 251485
rect 515711 251393 515745 251409
rect 515869 251469 515903 251485
rect 515869 251393 515903 251409
rect 515987 251469 516021 251485
rect 515987 251393 516021 251409
rect 516145 251469 516179 251485
rect 516145 251393 516179 251409
rect 516263 251469 516297 251485
rect 516263 251393 516297 251409
rect 516421 251469 516455 251485
rect 516421 251393 516455 251409
rect 516539 251469 516573 251485
rect 516539 251393 516573 251409
rect 516697 251469 516731 251485
rect 516697 251393 516731 251409
rect 516815 251469 516849 251485
rect 516815 251393 516849 251409
rect 516973 251469 517007 251485
rect 516973 251393 517007 251409
rect 517091 251469 517125 251485
rect 517091 251393 517125 251409
rect 517249 251469 517283 251485
rect 517249 251393 517283 251409
rect 503337 251325 503353 251359
rect 503421 251356 503437 251359
rect 503421 251325 503445 251356
rect 503613 251325 503629 251359
rect 503697 251325 503713 251359
rect 503889 251355 503905 251359
rect 503886 251325 503905 251355
rect 503973 251325 503989 251359
rect 504165 251351 504181 251359
rect 504162 251325 504181 251351
rect 504249 251325 504265 251359
rect 504441 251345 504457 251359
rect 504440 251325 504457 251345
rect 504525 251325 504541 251359
rect 504717 251341 504733 251359
rect 504716 251325 504733 251341
rect 504801 251325 504817 251359
rect 504993 251343 505009 251359
rect 504990 251325 505009 251343
rect 505077 251325 505093 251359
rect 505269 251341 505285 251359
rect 505268 251325 505285 251341
rect 505353 251325 505369 251359
rect 505545 251325 505561 251359
rect 505629 251325 505645 251359
rect 505821 251341 505837 251359
rect 505820 251325 505837 251341
rect 505905 251325 505921 251359
rect 506097 251325 506113 251359
rect 506181 251325 506197 251359
rect 506373 251351 506389 251359
rect 506370 251335 506389 251351
rect 506369 251325 506389 251335
rect 506457 251325 506473 251359
rect 506649 251351 506665 251359
rect 506646 251325 506665 251351
rect 506733 251325 506749 251359
rect 506925 251325 506941 251359
rect 507009 251325 507025 251359
rect 507201 251345 507217 251359
rect 507194 251325 507217 251345
rect 507285 251325 507301 251359
rect 507477 251325 507493 251359
rect 507561 251325 507577 251359
rect 507753 251345 507769 251359
rect 507752 251325 507769 251345
rect 507837 251325 507853 251359
rect 508029 251341 508045 251359
rect 508028 251325 508045 251341
rect 508113 251325 508129 251359
rect 508305 251349 508321 251359
rect 508302 251325 508321 251349
rect 508389 251325 508405 251359
rect 508581 251341 508597 251359
rect 508580 251325 508597 251341
rect 508665 251325 508681 251359
rect 508857 251343 508873 251359
rect 508850 251325 508873 251343
rect 508941 251325 508957 251359
rect 509133 251349 509149 251359
rect 509126 251325 509149 251349
rect 509217 251325 509233 251359
rect 509409 251355 509425 251359
rect 509408 251325 509425 251355
rect 509493 251325 509509 251359
rect 509685 251351 509701 251359
rect 509684 251325 509701 251351
rect 509769 251325 509785 251359
rect 509961 251351 509977 251359
rect 509958 251325 509977 251351
rect 510045 251325 510061 251359
rect 510237 251351 510253 251359
rect 510230 251325 510253 251351
rect 510321 251325 510337 251359
rect 510513 251351 510529 251359
rect 510512 251325 510529 251351
rect 510597 251325 510613 251359
rect 510789 251325 510805 251359
rect 510873 251325 510889 251359
rect 511065 251345 511081 251359
rect 511064 251325 511081 251345
rect 511149 251325 511165 251359
rect 511341 251325 511357 251359
rect 511425 251325 511441 251359
rect 511617 251325 511633 251359
rect 511701 251325 511717 251359
rect 511893 251337 511909 251359
rect 511886 251325 511909 251337
rect 511977 251325 511993 251359
rect 512169 251333 512185 251359
rect 512168 251325 512185 251333
rect 512253 251325 512269 251359
rect 512445 251325 512461 251359
rect 512529 251325 512545 251359
rect 512721 251333 512737 251359
rect 512720 251325 512737 251333
rect 512805 251325 512821 251359
rect 512997 251333 513013 251359
rect 512996 251325 513013 251333
rect 513081 251325 513097 251359
rect 513273 251349 513289 251359
rect 513266 251325 513289 251349
rect 513357 251325 513373 251359
rect 513549 251341 513565 251359
rect 513544 251325 513565 251341
rect 513633 251325 513649 251359
rect 513825 251325 513841 251359
rect 513909 251325 513925 251359
rect 514101 251325 514117 251359
rect 514185 251341 514201 251359
rect 514377 251345 514393 251359
rect 514185 251325 514206 251341
rect 503343 251116 503445 251325
rect 503614 251116 503712 251325
rect 503886 251116 503984 251325
rect 504162 251116 504260 251325
rect 504440 251116 504538 251325
rect 504716 251116 504814 251325
rect 504990 251116 505088 251325
rect 505268 251116 505366 251325
rect 505546 251116 505644 251325
rect 505820 251116 505918 251325
rect 506098 251116 506196 251325
rect 506369 251116 506469 251325
rect 506646 251116 506744 251325
rect 506926 251116 507024 251325
rect 507194 251116 507292 251325
rect 507478 251116 507576 251325
rect 507752 251116 507850 251325
rect 508028 251116 508126 251325
rect 508302 251116 508400 251325
rect 508580 251116 508678 251325
rect 508850 251116 508948 251325
rect 509126 251116 509224 251325
rect 509408 251116 509506 251325
rect 509684 251116 509782 251325
rect 509958 251310 510056 251325
rect 510230 251116 510328 251325
rect 510512 251116 510610 251325
rect 510790 251116 510888 251325
rect 511064 251116 511162 251325
rect 511342 251116 511440 251325
rect 511618 251116 511716 251325
rect 511886 251116 511984 251325
rect 512168 251116 512266 251325
rect 512446 251116 512544 251325
rect 512720 251116 512818 251325
rect 512996 251116 513094 251325
rect 513266 251116 513364 251325
rect 513544 251116 513642 251325
rect 513826 251116 513924 251325
rect 514108 251116 514206 251325
rect 514376 251325 514393 251345
rect 514461 251325 514477 251359
rect 514653 251345 514669 251359
rect 514652 251325 514669 251345
rect 514737 251325 514753 251359
rect 514929 251345 514945 251359
rect 514922 251325 514945 251345
rect 515013 251325 515029 251359
rect 515205 251351 515221 251359
rect 515200 251325 515221 251351
rect 515289 251325 515305 251359
rect 515481 251325 515497 251359
rect 515565 251325 515581 251359
rect 515757 251325 515773 251359
rect 515841 251351 515857 251359
rect 515841 251325 515860 251351
rect 516033 251349 516049 251359
rect 514376 251116 514474 251325
rect 514652 251116 514750 251325
rect 514922 251116 515020 251325
rect 515200 251116 515298 251325
rect 515482 251116 515580 251325
rect 515762 251116 515860 251325
rect 516028 251325 516049 251349
rect 516117 251325 516133 251359
rect 516309 251343 516325 251359
rect 516304 251325 516325 251343
rect 516393 251325 516409 251359
rect 516585 251349 516601 251359
rect 516584 251325 516601 251349
rect 516669 251325 516685 251359
rect 516861 251325 516877 251359
rect 516945 251349 516961 251359
rect 516945 251325 516966 251349
rect 517137 251325 517153 251359
rect 517221 251353 517237 251359
rect 517221 251325 517244 251353
rect 516028 251116 516126 251325
rect 516304 251116 516402 251325
rect 516584 251116 516682 251325
rect 516868 251116 516966 251325
rect 517146 251116 517244 251325
rect 517383 251267 517417 251283
rect 517735 251116 517833 251740
rect 413340 251085 427833 251116
rect 413340 251029 417346 251085
rect 417424 251029 427833 251085
rect 413340 251018 427833 251029
rect 503340 251085 517833 251116
rect 503340 251029 507346 251085
rect 507424 251029 517833 251085
rect 503340 251018 517833 251029
rect 322697 250489 337190 250520
rect 322697 250433 326703 250489
rect 326781 250433 337190 250489
rect 322697 250422 337190 250433
rect 239514 146062 239548 146078
rect 59497 146033 59531 146049
rect 59323 145993 59339 146027
rect 59373 145993 59389 146027
rect 59295 145934 59329 145950
rect 59295 145742 59329 145758
rect 59383 145934 59417 145950
rect 59383 145742 59417 145758
rect 59323 145665 59339 145699
rect 59373 145665 59389 145699
rect 239340 146022 239356 146056
rect 239390 146022 239406 146056
rect 239312 145972 239346 145988
rect 239312 145780 239346 145796
rect 239400 145972 239434 145988
rect 239400 145780 239434 145796
rect 239340 145712 239356 145746
rect 239390 145712 239406 145746
rect 509514 146062 509548 146078
rect 329497 146033 329531 146049
rect 329323 145993 329339 146027
rect 329373 145993 329389 146027
rect 329295 145934 329329 145950
rect 329295 145742 329329 145758
rect 329383 145934 329417 145950
rect 329383 145742 329417 145758
rect 239514 145690 239548 145706
rect 59497 145643 59531 145659
rect 149767 145665 149801 145681
rect 329323 145665 329339 145699
rect 329373 145665 329389 145699
rect 149521 145589 149537 145623
rect 149605 145589 149621 145623
rect 149475 145530 149509 145546
rect 149475 145338 149509 145354
rect 149633 145530 149667 145546
rect 149633 145338 149667 145354
rect 149521 145261 149537 145295
rect 149605 145261 149621 145295
rect 509340 146022 509356 146056
rect 509390 146022 509406 146056
rect 509312 145972 509346 145988
rect 509312 145780 509346 145796
rect 509400 145972 509434 145988
rect 509400 145780 509434 145796
rect 509340 145712 509356 145746
rect 509390 145712 509406 145746
rect 509514 145690 509548 145706
rect 329497 145643 329531 145659
rect 419767 145665 419801 145681
rect 419521 145589 419537 145623
rect 419605 145589 419621 145623
rect 419475 145530 419509 145546
rect 419475 145338 419509 145354
rect 419633 145530 419667 145546
rect 419633 145338 419667 145354
rect 419521 145261 419537 145295
rect 419605 145261 419621 145295
rect 149767 145203 149801 145219
rect 419767 145203 419801 145219
rect 149857 56097 149891 56113
rect 59514 56062 59548 56078
rect 59340 56022 59356 56056
rect 59390 56022 59406 56056
rect 59312 55972 59346 55988
rect 59312 55780 59346 55796
rect 59400 55972 59434 55988
rect 59400 55780 59434 55796
rect 59340 55712 59356 55746
rect 59390 55712 59406 55746
rect 149611 56021 149627 56055
rect 149695 56021 149711 56055
rect 149565 55971 149599 55987
rect 149565 55779 149599 55795
rect 149723 55971 149757 55987
rect 149723 55779 149757 55795
rect 149611 55711 149627 55745
rect 149695 55711 149711 55745
rect 59514 55690 59548 55706
rect 419857 56097 419891 56113
rect 329514 56062 329548 56078
rect 329340 56022 329356 56056
rect 329390 56022 329406 56056
rect 329312 55972 329346 55988
rect 239867 55807 239901 55823
rect 239621 55731 239637 55765
rect 239705 55731 239721 55765
rect 149857 55653 149891 55669
rect 239575 55681 239609 55697
rect 239575 55489 239609 55505
rect 239733 55681 239767 55697
rect 239733 55489 239767 55505
rect 239621 55421 239637 55455
rect 239705 55421 239721 55455
rect 329312 55780 329346 55796
rect 329400 55972 329434 55988
rect 329400 55780 329434 55796
rect 329340 55712 329356 55746
rect 329390 55712 329406 55746
rect 419611 56021 419627 56055
rect 419695 56021 419711 56055
rect 419565 55971 419599 55987
rect 419565 55779 419599 55795
rect 419723 55971 419757 55987
rect 419723 55779 419757 55795
rect 419611 55711 419627 55745
rect 419695 55711 419711 55745
rect 329514 55690 329548 55706
rect 509867 55807 509901 55823
rect 509621 55731 509637 55765
rect 509705 55731 509721 55765
rect 419857 55653 419891 55669
rect 509575 55681 509609 55697
rect 509575 55489 509609 55505
rect 509733 55681 509767 55697
rect 509733 55489 509767 55505
rect 509621 55421 509637 55455
rect 509705 55421 509721 55455
rect 239867 55363 239901 55379
rect 509867 55363 509901 55379
<< viali >>
rect 329158 657946 329192 657980
rect 329114 657720 329148 657896
rect 329202 657720 329236 657896
rect 329158 657636 329192 657670
rect 509158 657946 509192 657980
rect 509114 657720 509148 657896
rect 509202 657720 509236 657896
rect 509158 657636 509192 657670
rect 419339 657513 419407 657547
rect 419277 657278 419311 657454
rect 419435 657278 419469 657454
rect 419339 657185 419407 657219
rect 59627 656021 59695 656055
rect 59565 655795 59599 655971
rect 59723 655795 59757 655971
rect 59627 655711 59695 655745
rect 149356 656022 149390 656056
rect 149312 655796 149346 655972
rect 149400 655796 149434 655972
rect 149356 655712 149390 655746
rect 239339 655993 239373 656027
rect 239295 655758 239329 655934
rect 239383 655758 239417 655934
rect 239339 655665 239373 655699
rect 419429 582945 419497 582979
rect 419367 582719 419401 582895
rect 419525 582719 419559 582895
rect 419429 582635 419497 582669
rect 509439 582655 509507 582689
rect 509377 582429 509411 582605
rect 509535 582429 509569 582605
rect 509439 582345 509507 582379
rect 59627 581021 59695 581055
rect 59565 580795 59599 580971
rect 59723 580795 59757 580971
rect 59627 580711 59695 580745
rect 239356 581022 239390 581056
rect 149637 580731 149705 580765
rect 149575 580505 149609 580681
rect 149733 580505 149767 580681
rect 149637 580421 149705 580455
rect 239312 580796 239346 580972
rect 239400 580796 239434 580972
rect 239356 580712 239390 580746
rect 329537 580589 329605 580623
rect 329475 580354 329509 580530
rect 329633 580354 329667 580530
rect 329537 580261 329605 580295
rect 323904 492556 323958 492598
rect 323893 492197 323961 492231
rect 324169 492197 324237 492231
rect 324445 492197 324513 492231
rect 324721 492197 324789 492231
rect 324997 492197 325065 492231
rect 325273 492197 325341 492231
rect 325549 492197 325617 492231
rect 325825 492197 325893 492231
rect 326101 492197 326169 492231
rect 326377 492197 326445 492231
rect 326653 492197 326721 492231
rect 326929 492197 326997 492231
rect 327205 492197 327273 492231
rect 327481 492197 327549 492231
rect 327757 492197 327825 492231
rect 328033 492197 328101 492231
rect 328309 492197 328377 492231
rect 328585 492197 328653 492231
rect 328861 492197 328929 492231
rect 329137 492197 329205 492231
rect 329413 492197 329481 492231
rect 329689 492197 329757 492231
rect 329965 492197 330033 492231
rect 330241 492197 330309 492231
rect 330517 492197 330585 492231
rect 330793 492197 330861 492231
rect 331069 492197 331137 492231
rect 331345 492197 331413 492231
rect 331621 492197 331689 492231
rect 331897 492197 331965 492231
rect 332173 492197 332241 492231
rect 332449 492197 332517 492231
rect 332725 492197 332793 492231
rect 333001 492197 333069 492231
rect 333277 492197 333345 492231
rect 333553 492197 333621 492231
rect 333829 492197 333897 492231
rect 334105 492197 334173 492231
rect 334381 492197 334449 492231
rect 334657 492197 334725 492231
rect 334933 492197 335001 492231
rect 335209 492197 335277 492231
rect 335485 492197 335553 492231
rect 335761 492197 335829 492231
rect 336037 492197 336105 492231
rect 336313 492197 336381 492231
rect 336589 492197 336657 492231
rect 336865 492197 336933 492231
rect 337141 492197 337209 492231
rect 337417 492197 337485 492231
rect 337693 492197 337761 492231
rect 323831 492087 323865 492147
rect 323989 492087 324023 492147
rect 324107 492087 324141 492147
rect 324265 492087 324299 492147
rect 324383 492087 324417 492147
rect 324541 492087 324575 492147
rect 324659 492087 324693 492147
rect 324817 492087 324851 492147
rect 324935 492087 324969 492147
rect 325093 492087 325127 492147
rect 325211 492087 325245 492147
rect 325369 492087 325403 492147
rect 325487 492087 325521 492147
rect 325645 492087 325679 492147
rect 325763 492087 325797 492147
rect 325921 492087 325955 492147
rect 326039 492087 326073 492147
rect 326197 492087 326231 492147
rect 326315 492087 326349 492147
rect 326473 492087 326507 492147
rect 326591 492087 326625 492147
rect 326749 492087 326783 492147
rect 326867 492087 326901 492147
rect 327025 492087 327059 492147
rect 327143 492087 327177 492147
rect 327301 492087 327335 492147
rect 327419 492087 327453 492147
rect 327577 492087 327611 492147
rect 327695 492087 327729 492147
rect 327853 492087 327887 492147
rect 327971 492087 328005 492147
rect 328129 492087 328163 492147
rect 328247 492087 328281 492147
rect 328405 492087 328439 492147
rect 328523 492087 328557 492147
rect 328681 492087 328715 492147
rect 328799 492087 328833 492147
rect 328957 492087 328991 492147
rect 329075 492087 329109 492147
rect 329233 492087 329267 492147
rect 329351 492087 329385 492147
rect 329509 492087 329543 492147
rect 329627 492087 329661 492147
rect 329785 492087 329819 492147
rect 329903 492087 329937 492147
rect 330061 492087 330095 492147
rect 330179 492087 330213 492147
rect 330337 492087 330371 492147
rect 330455 492087 330489 492147
rect 330613 492087 330647 492147
rect 330731 492087 330765 492147
rect 330889 492087 330923 492147
rect 331007 492087 331041 492147
rect 331165 492087 331199 492147
rect 331283 492087 331317 492147
rect 331441 492087 331475 492147
rect 331559 492087 331593 492147
rect 331717 492087 331751 492147
rect 331835 492087 331869 492147
rect 331993 492087 332027 492147
rect 332111 492087 332145 492147
rect 332269 492087 332303 492147
rect 332387 492087 332421 492147
rect 332545 492087 332579 492147
rect 332663 492087 332697 492147
rect 332821 492087 332855 492147
rect 332939 492087 332973 492147
rect 333097 492087 333131 492147
rect 333215 492087 333249 492147
rect 333373 492087 333407 492147
rect 333491 492087 333525 492147
rect 333649 492087 333683 492147
rect 333767 492087 333801 492147
rect 333925 492087 333959 492147
rect 334043 492087 334077 492147
rect 334201 492087 334235 492147
rect 334319 492087 334353 492147
rect 334477 492087 334511 492147
rect 334595 492087 334629 492147
rect 334753 492087 334787 492147
rect 334871 492087 334905 492147
rect 335029 492087 335063 492147
rect 335147 492087 335181 492147
rect 335305 492087 335339 492147
rect 335423 492087 335457 492147
rect 335581 492087 335615 492147
rect 335699 492087 335733 492147
rect 335857 492087 335891 492147
rect 335975 492087 336009 492147
rect 336133 492087 336167 492147
rect 336251 492087 336285 492147
rect 336409 492087 336443 492147
rect 336527 492087 336561 492147
rect 336685 492087 336719 492147
rect 336803 492087 336837 492147
rect 336961 492087 336995 492147
rect 337079 492087 337113 492147
rect 337237 492087 337271 492147
rect 337355 492087 337389 492147
rect 337513 492087 337547 492147
rect 337631 492087 337665 492147
rect 337789 492087 337823 492147
rect 323893 492003 323961 492037
rect 324169 492003 324237 492037
rect 324445 492003 324513 492037
rect 324721 492003 324789 492037
rect 324997 492003 325065 492037
rect 325273 492003 325341 492037
rect 325549 492003 325617 492037
rect 325825 492003 325893 492037
rect 326101 492003 326169 492037
rect 326377 492003 326445 492037
rect 326653 492003 326721 492037
rect 326929 492003 326997 492037
rect 327205 492003 327273 492037
rect 327481 492003 327549 492037
rect 327757 492003 327825 492037
rect 328033 492003 328101 492037
rect 328309 492003 328377 492037
rect 328585 492003 328653 492037
rect 328861 492003 328929 492037
rect 329137 492003 329205 492037
rect 329413 492003 329481 492037
rect 329689 492003 329757 492037
rect 329965 492003 330033 492037
rect 330241 492003 330309 492037
rect 330517 492003 330585 492037
rect 330793 492003 330861 492037
rect 331069 492003 331137 492037
rect 331345 492003 331413 492037
rect 331621 492003 331689 492037
rect 331897 492003 331965 492037
rect 332173 492003 332241 492037
rect 332449 492003 332517 492037
rect 332725 492003 332793 492037
rect 333001 492003 333069 492037
rect 333277 492003 333345 492037
rect 333553 492003 333621 492037
rect 333829 492003 333897 492037
rect 334105 492003 334173 492037
rect 334381 492003 334449 492037
rect 334657 492003 334725 492037
rect 58903 491809 58971 491843
rect 59179 491809 59247 491843
rect 59455 491809 59523 491843
rect 59731 491809 59799 491843
rect 60007 491809 60075 491843
rect 60283 491809 60351 491843
rect 60559 491809 60627 491843
rect 60835 491809 60903 491843
rect 61111 491809 61179 491843
rect 61387 491809 61455 491843
rect 58841 491699 58875 491759
rect 58999 491699 59033 491759
rect 59117 491699 59151 491759
rect 59275 491699 59309 491759
rect 59393 491699 59427 491759
rect 59551 491699 59585 491759
rect 59669 491699 59703 491759
rect 59827 491699 59861 491759
rect 59945 491699 59979 491759
rect 60103 491699 60137 491759
rect 60221 491699 60255 491759
rect 60379 491699 60413 491759
rect 60497 491699 60531 491759
rect 60655 491699 60689 491759
rect 60773 491699 60807 491759
rect 60931 491699 60965 491759
rect 61049 491699 61083 491759
rect 61207 491699 61241 491759
rect 61325 491699 61359 491759
rect 61483 491699 61517 491759
rect 58903 491615 58971 491649
rect 59179 491615 59247 491649
rect 59455 491615 59523 491649
rect 59731 491615 59799 491649
rect 60007 491615 60075 491649
rect 60283 491615 60351 491649
rect 60559 491615 60627 491649
rect 60835 491615 60903 491649
rect 61111 491615 61179 491649
rect 61387 491615 61455 491649
rect 143353 491519 143421 491553
rect 143629 491519 143697 491553
rect 143905 491519 143973 491553
rect 144181 491519 144249 491553
rect 144457 491519 144525 491553
rect 144733 491519 144801 491553
rect 145009 491519 145077 491553
rect 145285 491519 145353 491553
rect 145561 491519 145629 491553
rect 145837 491519 145905 491553
rect 146113 491519 146181 491553
rect 146389 491519 146457 491553
rect 146665 491519 146733 491553
rect 146941 491519 147009 491553
rect 147217 491519 147285 491553
rect 147493 491519 147561 491553
rect 147769 491519 147837 491553
rect 148045 491519 148113 491553
rect 148321 491519 148389 491553
rect 148597 491519 148665 491553
rect 148873 491519 148941 491553
rect 149149 491519 149217 491553
rect 149425 491519 149493 491553
rect 149701 491519 149769 491553
rect 149977 491519 150045 491553
rect 150253 491519 150321 491553
rect 150529 491519 150597 491553
rect 150805 491519 150873 491553
rect 151081 491519 151149 491553
rect 151357 491519 151425 491553
rect 151633 491519 151701 491553
rect 151909 491519 151977 491553
rect 152185 491519 152253 491553
rect 152461 491519 152529 491553
rect 152737 491519 152805 491553
rect 153013 491519 153081 491553
rect 153289 491519 153357 491553
rect 153565 491519 153633 491553
rect 153841 491519 153909 491553
rect 154117 491519 154185 491553
rect 154393 491519 154461 491553
rect 154669 491519 154737 491553
rect 154945 491519 155013 491553
rect 155221 491519 155289 491553
rect 155497 491519 155565 491553
rect 155773 491519 155841 491553
rect 156049 491519 156117 491553
rect 156325 491519 156393 491553
rect 156601 491519 156669 491553
rect 156877 491519 156945 491553
rect 157153 491519 157221 491553
rect 143291 491409 143325 491469
rect 143449 491409 143483 491469
rect 143567 491409 143601 491469
rect 143725 491409 143759 491469
rect 143843 491409 143877 491469
rect 144001 491409 144035 491469
rect 144119 491409 144153 491469
rect 144277 491409 144311 491469
rect 144395 491409 144429 491469
rect 144553 491409 144587 491469
rect 144671 491409 144705 491469
rect 144829 491409 144863 491469
rect 144947 491409 144981 491469
rect 145105 491409 145139 491469
rect 145223 491409 145257 491469
rect 145381 491409 145415 491469
rect 145499 491409 145533 491469
rect 145657 491409 145691 491469
rect 145775 491409 145809 491469
rect 145933 491409 145967 491469
rect 146051 491409 146085 491469
rect 146209 491409 146243 491469
rect 146327 491409 146361 491469
rect 146485 491409 146519 491469
rect 146603 491409 146637 491469
rect 146761 491409 146795 491469
rect 146879 491409 146913 491469
rect 147037 491409 147071 491469
rect 147155 491409 147189 491469
rect 147313 491409 147347 491469
rect 147431 491409 147465 491469
rect 147589 491409 147623 491469
rect 147707 491409 147741 491469
rect 147865 491409 147899 491469
rect 147983 491409 148017 491469
rect 148141 491409 148175 491469
rect 148259 491409 148293 491469
rect 148417 491409 148451 491469
rect 148535 491409 148569 491469
rect 148693 491409 148727 491469
rect 148811 491409 148845 491469
rect 148969 491409 149003 491469
rect 149087 491409 149121 491469
rect 149245 491409 149279 491469
rect 149363 491409 149397 491469
rect 149521 491409 149555 491469
rect 149639 491409 149673 491469
rect 149797 491409 149831 491469
rect 149915 491409 149949 491469
rect 150073 491409 150107 491469
rect 150191 491409 150225 491469
rect 150349 491409 150383 491469
rect 150467 491409 150501 491469
rect 150625 491409 150659 491469
rect 150743 491409 150777 491469
rect 150901 491409 150935 491469
rect 151019 491409 151053 491469
rect 151177 491409 151211 491469
rect 151295 491409 151329 491469
rect 151453 491409 151487 491469
rect 151571 491409 151605 491469
rect 151729 491409 151763 491469
rect 151847 491409 151881 491469
rect 152005 491409 152039 491469
rect 152123 491409 152157 491469
rect 152281 491409 152315 491469
rect 152399 491409 152433 491469
rect 152557 491409 152591 491469
rect 152675 491409 152709 491469
rect 152833 491409 152867 491469
rect 152951 491409 152985 491469
rect 153109 491409 153143 491469
rect 153227 491409 153261 491469
rect 153385 491409 153419 491469
rect 153503 491409 153537 491469
rect 153661 491409 153695 491469
rect 153779 491409 153813 491469
rect 153937 491409 153971 491469
rect 154055 491409 154089 491469
rect 154213 491409 154247 491469
rect 154331 491409 154365 491469
rect 154489 491409 154523 491469
rect 154607 491409 154641 491469
rect 154765 491409 154799 491469
rect 154883 491409 154917 491469
rect 155041 491409 155075 491469
rect 155159 491409 155193 491469
rect 155317 491409 155351 491469
rect 155435 491409 155469 491469
rect 155593 491409 155627 491469
rect 155711 491409 155745 491469
rect 155869 491409 155903 491469
rect 155987 491409 156021 491469
rect 156145 491409 156179 491469
rect 156263 491409 156297 491469
rect 156421 491409 156455 491469
rect 156539 491409 156573 491469
rect 156697 491409 156731 491469
rect 156815 491409 156849 491469
rect 156973 491409 157007 491469
rect 157091 491409 157125 491469
rect 157249 491409 157283 491469
rect 59566 491290 59638 491334
rect 143353 491325 143421 491359
rect 143629 491325 143697 491359
rect 143905 491325 143973 491359
rect 144181 491325 144249 491359
rect 144457 491325 144525 491359
rect 144733 491325 144801 491359
rect 145009 491325 145077 491359
rect 145285 491325 145353 491359
rect 145561 491325 145629 491359
rect 145837 491325 145905 491359
rect 146113 491325 146181 491359
rect 146389 491325 146457 491359
rect 146665 491325 146733 491359
rect 146941 491325 147009 491359
rect 147217 491325 147285 491359
rect 147493 491325 147561 491359
rect 147769 491325 147837 491359
rect 148045 491325 148113 491359
rect 148321 491325 148389 491359
rect 148597 491325 148665 491359
rect 148873 491325 148941 491359
rect 149149 491325 149217 491359
rect 149425 491325 149493 491359
rect 149701 491325 149769 491359
rect 149977 491325 150045 491359
rect 150253 491325 150321 491359
rect 150529 491325 150597 491359
rect 150805 491325 150873 491359
rect 151081 491325 151149 491359
rect 151357 491325 151425 491359
rect 151633 491325 151701 491359
rect 151909 491325 151977 491359
rect 152185 491325 152253 491359
rect 152461 491325 152529 491359
rect 152737 491325 152805 491359
rect 153013 491325 153081 491359
rect 153289 491325 153357 491359
rect 153565 491325 153633 491359
rect 153841 491325 153909 491359
rect 154117 491325 154185 491359
rect 154393 491325 154461 491359
rect 154669 491325 154737 491359
rect 154945 491325 155013 491359
rect 155221 491325 155289 491359
rect 155497 491325 155565 491359
rect 155773 491325 155841 491359
rect 156049 491325 156117 491359
rect 156325 491325 156393 491359
rect 156601 491325 156669 491359
rect 156877 491325 156945 491359
rect 157153 491325 157221 491359
rect 334933 492003 335001 492037
rect 335209 492003 335277 492037
rect 335485 492003 335553 492037
rect 335761 492003 335829 492037
rect 336037 492003 336105 492037
rect 336313 492003 336381 492037
rect 336589 492003 336657 492037
rect 336865 492003 336933 492037
rect 337141 492003 337209 492037
rect 337417 492003 337485 492037
rect 337693 492003 337761 492037
rect 327886 491706 327964 491762
rect 323904 491644 323958 491686
rect 418902 491481 418970 491515
rect 419178 491481 419246 491515
rect 419454 491481 419522 491515
rect 419730 491481 419798 491515
rect 420006 491481 420074 491515
rect 418840 491371 418874 491431
rect 418998 491371 419032 491431
rect 419116 491371 419150 491431
rect 419274 491371 419308 491431
rect 419392 491371 419426 491431
rect 419550 491371 419584 491431
rect 419668 491371 419702 491431
rect 419826 491371 419860 491431
rect 419944 491371 419978 491431
rect 420102 491371 420136 491431
rect 418902 491287 418970 491321
rect 419178 491287 419246 491321
rect 419454 491287 419522 491321
rect 419730 491287 419798 491321
rect 420006 491287 420074 491321
rect 418923 491210 418961 491244
rect 508903 491809 508971 491843
rect 509179 491809 509247 491843
rect 509455 491809 509523 491843
rect 509731 491809 509799 491843
rect 510007 491809 510075 491843
rect 510283 491809 510351 491843
rect 510559 491809 510627 491843
rect 510835 491809 510903 491843
rect 511111 491809 511179 491843
rect 511387 491809 511455 491843
rect 508841 491699 508875 491759
rect 508999 491699 509033 491759
rect 509117 491699 509151 491759
rect 509275 491699 509309 491759
rect 509393 491699 509427 491759
rect 509551 491699 509585 491759
rect 509669 491699 509703 491759
rect 509827 491699 509861 491759
rect 509945 491699 509979 491759
rect 510103 491699 510137 491759
rect 510221 491699 510255 491759
rect 510379 491699 510413 491759
rect 510497 491699 510531 491759
rect 510655 491699 510689 491759
rect 510773 491699 510807 491759
rect 510931 491699 510965 491759
rect 511049 491699 511083 491759
rect 511207 491699 511241 491759
rect 511325 491699 511359 491759
rect 511483 491699 511517 491759
rect 508903 491615 508971 491649
rect 509179 491615 509247 491649
rect 509455 491615 509523 491649
rect 509731 491615 509799 491649
rect 510007 491615 510075 491649
rect 510283 491615 510351 491649
rect 510559 491615 510627 491649
rect 510835 491615 510903 491649
rect 511111 491615 511179 491649
rect 511387 491615 511455 491649
rect 509566 491290 509638 491334
rect 147346 491029 147424 491085
rect 232710 490923 232778 490957
rect 232986 490923 233054 490957
rect 233262 490923 233330 490957
rect 233538 490923 233606 490957
rect 233814 490923 233882 490957
rect 234090 490923 234158 490957
rect 234366 490923 234434 490957
rect 234642 490923 234710 490957
rect 234918 490923 234986 490957
rect 235194 490923 235262 490957
rect 235470 490923 235538 490957
rect 235746 490923 235814 490957
rect 236022 490923 236090 490957
rect 236298 490923 236366 490957
rect 236574 490923 236642 490957
rect 236850 490923 236918 490957
rect 237126 490923 237194 490957
rect 237402 490923 237470 490957
rect 237678 490923 237746 490957
rect 237954 490923 238022 490957
rect 238230 490923 238298 490957
rect 238506 490923 238574 490957
rect 238782 490923 238850 490957
rect 239058 490923 239126 490957
rect 239334 490923 239402 490957
rect 239610 490923 239678 490957
rect 239886 490923 239954 490957
rect 240162 490923 240230 490957
rect 240438 490923 240506 490957
rect 240714 490923 240782 490957
rect 240990 490923 241058 490957
rect 241266 490923 241334 490957
rect 241542 490923 241610 490957
rect 241818 490923 241886 490957
rect 242094 490923 242162 490957
rect 242370 490923 242438 490957
rect 242646 490923 242714 490957
rect 242922 490923 242990 490957
rect 243198 490923 243266 490957
rect 243474 490923 243542 490957
rect 243750 490923 243818 490957
rect 244026 490923 244094 490957
rect 244302 490923 244370 490957
rect 244578 490923 244646 490957
rect 244854 490923 244922 490957
rect 245130 490923 245198 490957
rect 245406 490923 245474 490957
rect 245682 490923 245750 490957
rect 245958 490923 246026 490957
rect 246234 490923 246302 490957
rect 246510 490923 246578 490957
rect 232648 490813 232682 490873
rect 232806 490813 232840 490873
rect 232924 490813 232958 490873
rect 233082 490813 233116 490873
rect 233200 490813 233234 490873
rect 233358 490813 233392 490873
rect 233476 490813 233510 490873
rect 233634 490813 233668 490873
rect 233752 490813 233786 490873
rect 233910 490813 233944 490873
rect 234028 490813 234062 490873
rect 234186 490813 234220 490873
rect 234304 490813 234338 490873
rect 234462 490813 234496 490873
rect 234580 490813 234614 490873
rect 234738 490813 234772 490873
rect 234856 490813 234890 490873
rect 235014 490813 235048 490873
rect 235132 490813 235166 490873
rect 235290 490813 235324 490873
rect 235408 490813 235442 490873
rect 235566 490813 235600 490873
rect 235684 490813 235718 490873
rect 235842 490813 235876 490873
rect 235960 490813 235994 490873
rect 236118 490813 236152 490873
rect 236236 490813 236270 490873
rect 236394 490813 236428 490873
rect 236512 490813 236546 490873
rect 236670 490813 236704 490873
rect 236788 490813 236822 490873
rect 236946 490813 236980 490873
rect 237064 490813 237098 490873
rect 237222 490813 237256 490873
rect 237340 490813 237374 490873
rect 237498 490813 237532 490873
rect 237616 490813 237650 490873
rect 237774 490813 237808 490873
rect 237892 490813 237926 490873
rect 238050 490813 238084 490873
rect 238168 490813 238202 490873
rect 238326 490813 238360 490873
rect 238444 490813 238478 490873
rect 238602 490813 238636 490873
rect 238720 490813 238754 490873
rect 238878 490813 238912 490873
rect 238996 490813 239030 490873
rect 239154 490813 239188 490873
rect 239272 490813 239306 490873
rect 239430 490813 239464 490873
rect 239548 490813 239582 490873
rect 239706 490813 239740 490873
rect 239824 490813 239858 490873
rect 239982 490813 240016 490873
rect 240100 490813 240134 490873
rect 240258 490813 240292 490873
rect 240376 490813 240410 490873
rect 240534 490813 240568 490873
rect 240652 490813 240686 490873
rect 240810 490813 240844 490873
rect 240928 490813 240962 490873
rect 241086 490813 241120 490873
rect 241204 490813 241238 490873
rect 241362 490813 241396 490873
rect 241480 490813 241514 490873
rect 241638 490813 241672 490873
rect 241756 490813 241790 490873
rect 241914 490813 241948 490873
rect 242032 490813 242066 490873
rect 242190 490813 242224 490873
rect 242308 490813 242342 490873
rect 242466 490813 242500 490873
rect 242584 490813 242618 490873
rect 242742 490813 242776 490873
rect 242860 490813 242894 490873
rect 243018 490813 243052 490873
rect 243136 490813 243170 490873
rect 243294 490813 243328 490873
rect 243412 490813 243446 490873
rect 243570 490813 243604 490873
rect 243688 490813 243722 490873
rect 243846 490813 243880 490873
rect 243964 490813 243998 490873
rect 244122 490813 244156 490873
rect 244240 490813 244274 490873
rect 244398 490813 244432 490873
rect 244516 490813 244550 490873
rect 244674 490813 244708 490873
rect 244792 490813 244826 490873
rect 244950 490813 244984 490873
rect 245068 490813 245102 490873
rect 245226 490813 245260 490873
rect 245344 490813 245378 490873
rect 245502 490813 245536 490873
rect 245620 490813 245654 490873
rect 245778 490813 245812 490873
rect 245896 490813 245930 490873
rect 246054 490813 246088 490873
rect 246172 490813 246206 490873
rect 246330 490813 246364 490873
rect 246448 490813 246482 490873
rect 246606 490813 246640 490873
rect 232710 490729 232778 490763
rect 232986 490729 233054 490763
rect 233262 490729 233330 490763
rect 233538 490729 233606 490763
rect 233814 490729 233882 490763
rect 234090 490729 234158 490763
rect 234366 490729 234434 490763
rect 234642 490729 234710 490763
rect 234918 490729 234986 490763
rect 235194 490729 235262 490763
rect 235470 490729 235538 490763
rect 235746 490729 235814 490763
rect 236022 490729 236090 490763
rect 236298 490729 236366 490763
rect 236574 490729 236642 490763
rect 236850 490729 236918 490763
rect 237126 490729 237194 490763
rect 237402 490729 237470 490763
rect 237678 490729 237746 490763
rect 237954 490729 238022 490763
rect 238230 490729 238298 490763
rect 238506 490729 238574 490763
rect 238782 490729 238850 490763
rect 239058 490729 239126 490763
rect 239334 490729 239402 490763
rect 239610 490729 239678 490763
rect 239886 490729 239954 490763
rect 240162 490729 240230 490763
rect 240438 490729 240506 490763
rect 240714 490729 240782 490763
rect 240990 490729 241058 490763
rect 241266 490729 241334 490763
rect 241542 490729 241610 490763
rect 241818 490729 241886 490763
rect 242094 490729 242162 490763
rect 242370 490729 242438 490763
rect 242646 490729 242714 490763
rect 242922 490729 242990 490763
rect 243198 490729 243266 490763
rect 243474 490729 243542 490763
rect 243750 490729 243818 490763
rect 244026 490729 244094 490763
rect 244302 490729 244370 490763
rect 244578 490729 244646 490763
rect 244854 490729 244922 490763
rect 245130 490729 245198 490763
rect 245406 490729 245474 490763
rect 245682 490729 245750 490763
rect 245958 490729 246026 490763
rect 246234 490729 246302 490763
rect 246510 490729 246578 490763
rect 236703 490433 236781 490489
rect 323904 372556 323958 372598
rect 323893 372197 323961 372231
rect 324169 372197 324237 372231
rect 324445 372197 324513 372231
rect 324721 372197 324789 372231
rect 324997 372197 325065 372231
rect 325273 372197 325341 372231
rect 325549 372197 325617 372231
rect 325825 372197 325893 372231
rect 326101 372197 326169 372231
rect 326377 372197 326445 372231
rect 326653 372197 326721 372231
rect 326929 372197 326997 372231
rect 327205 372197 327273 372231
rect 327481 372197 327549 372231
rect 327757 372197 327825 372231
rect 328033 372197 328101 372231
rect 328309 372197 328377 372231
rect 328585 372197 328653 372231
rect 328861 372197 328929 372231
rect 329137 372197 329205 372231
rect 329413 372197 329481 372231
rect 329689 372197 329757 372231
rect 329965 372197 330033 372231
rect 330241 372197 330309 372231
rect 330517 372197 330585 372231
rect 330793 372197 330861 372231
rect 331069 372197 331137 372231
rect 331345 372197 331413 372231
rect 331621 372197 331689 372231
rect 331897 372197 331965 372231
rect 332173 372197 332241 372231
rect 332449 372197 332517 372231
rect 332725 372197 332793 372231
rect 333001 372197 333069 372231
rect 333277 372197 333345 372231
rect 333553 372197 333621 372231
rect 333829 372197 333897 372231
rect 334105 372197 334173 372231
rect 334381 372197 334449 372231
rect 334657 372197 334725 372231
rect 334933 372197 335001 372231
rect 335209 372197 335277 372231
rect 335485 372197 335553 372231
rect 335761 372197 335829 372231
rect 336037 372197 336105 372231
rect 336313 372197 336381 372231
rect 336589 372197 336657 372231
rect 336865 372197 336933 372231
rect 337141 372197 337209 372231
rect 337417 372197 337485 372231
rect 337693 372197 337761 372231
rect 323831 372087 323865 372147
rect 323989 372087 324023 372147
rect 324107 372087 324141 372147
rect 324265 372087 324299 372147
rect 324383 372087 324417 372147
rect 324541 372087 324575 372147
rect 324659 372087 324693 372147
rect 324817 372087 324851 372147
rect 324935 372087 324969 372147
rect 325093 372087 325127 372147
rect 325211 372087 325245 372147
rect 325369 372087 325403 372147
rect 325487 372087 325521 372147
rect 325645 372087 325679 372147
rect 325763 372087 325797 372147
rect 325921 372087 325955 372147
rect 326039 372087 326073 372147
rect 326197 372087 326231 372147
rect 326315 372087 326349 372147
rect 326473 372087 326507 372147
rect 326591 372087 326625 372147
rect 326749 372087 326783 372147
rect 326867 372087 326901 372147
rect 327025 372087 327059 372147
rect 327143 372087 327177 372147
rect 327301 372087 327335 372147
rect 327419 372087 327453 372147
rect 327577 372087 327611 372147
rect 327695 372087 327729 372147
rect 327853 372087 327887 372147
rect 327971 372087 328005 372147
rect 328129 372087 328163 372147
rect 328247 372087 328281 372147
rect 328405 372087 328439 372147
rect 328523 372087 328557 372147
rect 328681 372087 328715 372147
rect 328799 372087 328833 372147
rect 328957 372087 328991 372147
rect 329075 372087 329109 372147
rect 329233 372087 329267 372147
rect 329351 372087 329385 372147
rect 329509 372087 329543 372147
rect 329627 372087 329661 372147
rect 329785 372087 329819 372147
rect 329903 372087 329937 372147
rect 330061 372087 330095 372147
rect 330179 372087 330213 372147
rect 330337 372087 330371 372147
rect 330455 372087 330489 372147
rect 330613 372087 330647 372147
rect 330731 372087 330765 372147
rect 330889 372087 330923 372147
rect 331007 372087 331041 372147
rect 331165 372087 331199 372147
rect 331283 372087 331317 372147
rect 331441 372087 331475 372147
rect 331559 372087 331593 372147
rect 331717 372087 331751 372147
rect 331835 372087 331869 372147
rect 331993 372087 332027 372147
rect 332111 372087 332145 372147
rect 332269 372087 332303 372147
rect 332387 372087 332421 372147
rect 332545 372087 332579 372147
rect 332663 372087 332697 372147
rect 332821 372087 332855 372147
rect 332939 372087 332973 372147
rect 333097 372087 333131 372147
rect 333215 372087 333249 372147
rect 333373 372087 333407 372147
rect 333491 372087 333525 372147
rect 333649 372087 333683 372147
rect 333767 372087 333801 372147
rect 333925 372087 333959 372147
rect 334043 372087 334077 372147
rect 334201 372087 334235 372147
rect 334319 372087 334353 372147
rect 334477 372087 334511 372147
rect 334595 372087 334629 372147
rect 334753 372087 334787 372147
rect 334871 372087 334905 372147
rect 335029 372087 335063 372147
rect 335147 372087 335181 372147
rect 335305 372087 335339 372147
rect 335423 372087 335457 372147
rect 335581 372087 335615 372147
rect 335699 372087 335733 372147
rect 335857 372087 335891 372147
rect 335975 372087 336009 372147
rect 336133 372087 336167 372147
rect 336251 372087 336285 372147
rect 336409 372087 336443 372147
rect 336527 372087 336561 372147
rect 336685 372087 336719 372147
rect 336803 372087 336837 372147
rect 336961 372087 336995 372147
rect 337079 372087 337113 372147
rect 337237 372087 337271 372147
rect 337355 372087 337389 372147
rect 337513 372087 337547 372147
rect 337631 372087 337665 372147
rect 337789 372087 337823 372147
rect 323893 372003 323961 372037
rect 324169 372003 324237 372037
rect 324445 372003 324513 372037
rect 324721 372003 324789 372037
rect 324997 372003 325065 372037
rect 325273 372003 325341 372037
rect 325549 372003 325617 372037
rect 325825 372003 325893 372037
rect 326101 372003 326169 372037
rect 326377 372003 326445 372037
rect 326653 372003 326721 372037
rect 326929 372003 326997 372037
rect 327205 372003 327273 372037
rect 327481 372003 327549 372037
rect 327757 372003 327825 372037
rect 328033 372003 328101 372037
rect 328309 372003 328377 372037
rect 328585 372003 328653 372037
rect 328861 372003 328929 372037
rect 329137 372003 329205 372037
rect 329413 372003 329481 372037
rect 329689 372003 329757 372037
rect 329965 372003 330033 372037
rect 330241 372003 330309 372037
rect 330517 372003 330585 372037
rect 330793 372003 330861 372037
rect 331069 372003 331137 372037
rect 331345 372003 331413 372037
rect 331621 372003 331689 372037
rect 331897 372003 331965 372037
rect 332173 372003 332241 372037
rect 332449 372003 332517 372037
rect 332725 372003 332793 372037
rect 333001 372003 333069 372037
rect 333277 372003 333345 372037
rect 333553 372003 333621 372037
rect 333829 372003 333897 372037
rect 334105 372003 334173 372037
rect 334381 372003 334449 372037
rect 334657 372003 334725 372037
rect 53353 371519 53421 371553
rect 53629 371519 53697 371553
rect 53905 371519 53973 371553
rect 54181 371519 54249 371553
rect 54457 371519 54525 371553
rect 54733 371519 54801 371553
rect 55009 371519 55077 371553
rect 55285 371519 55353 371553
rect 55561 371519 55629 371553
rect 55837 371519 55905 371553
rect 56113 371519 56181 371553
rect 56389 371519 56457 371553
rect 56665 371519 56733 371553
rect 56941 371519 57009 371553
rect 57217 371519 57285 371553
rect 57493 371519 57561 371553
rect 57769 371519 57837 371553
rect 58045 371519 58113 371553
rect 58321 371519 58389 371553
rect 58597 371519 58665 371553
rect 58873 371519 58941 371553
rect 59149 371519 59217 371553
rect 59425 371519 59493 371553
rect 59701 371519 59769 371553
rect 59977 371519 60045 371553
rect 60253 371519 60321 371553
rect 60529 371519 60597 371553
rect 60805 371519 60873 371553
rect 61081 371519 61149 371553
rect 61357 371519 61425 371553
rect 61633 371519 61701 371553
rect 61909 371519 61977 371553
rect 62185 371519 62253 371553
rect 62461 371519 62529 371553
rect 62737 371519 62805 371553
rect 63013 371519 63081 371553
rect 63289 371519 63357 371553
rect 63565 371519 63633 371553
rect 63841 371519 63909 371553
rect 64117 371519 64185 371553
rect 64393 371519 64461 371553
rect 64669 371519 64737 371553
rect 64945 371519 65013 371553
rect 65221 371519 65289 371553
rect 65497 371519 65565 371553
rect 65773 371519 65841 371553
rect 66049 371519 66117 371553
rect 66325 371519 66393 371553
rect 66601 371519 66669 371553
rect 66877 371519 66945 371553
rect 67153 371519 67221 371553
rect 53291 371409 53325 371469
rect 53449 371409 53483 371469
rect 53567 371409 53601 371469
rect 53725 371409 53759 371469
rect 53843 371409 53877 371469
rect 54001 371409 54035 371469
rect 54119 371409 54153 371469
rect 54277 371409 54311 371469
rect 54395 371409 54429 371469
rect 54553 371409 54587 371469
rect 54671 371409 54705 371469
rect 54829 371409 54863 371469
rect 54947 371409 54981 371469
rect 55105 371409 55139 371469
rect 55223 371409 55257 371469
rect 55381 371409 55415 371469
rect 55499 371409 55533 371469
rect 55657 371409 55691 371469
rect 55775 371409 55809 371469
rect 55933 371409 55967 371469
rect 56051 371409 56085 371469
rect 56209 371409 56243 371469
rect 56327 371409 56361 371469
rect 56485 371409 56519 371469
rect 56603 371409 56637 371469
rect 56761 371409 56795 371469
rect 56879 371409 56913 371469
rect 57037 371409 57071 371469
rect 57155 371409 57189 371469
rect 57313 371409 57347 371469
rect 57431 371409 57465 371469
rect 57589 371409 57623 371469
rect 57707 371409 57741 371469
rect 57865 371409 57899 371469
rect 57983 371409 58017 371469
rect 58141 371409 58175 371469
rect 58259 371409 58293 371469
rect 58417 371409 58451 371469
rect 58535 371409 58569 371469
rect 58693 371409 58727 371469
rect 58811 371409 58845 371469
rect 58969 371409 59003 371469
rect 59087 371409 59121 371469
rect 59245 371409 59279 371469
rect 59363 371409 59397 371469
rect 59521 371409 59555 371469
rect 59639 371409 59673 371469
rect 59797 371409 59831 371469
rect 59915 371409 59949 371469
rect 60073 371409 60107 371469
rect 60191 371409 60225 371469
rect 60349 371409 60383 371469
rect 60467 371409 60501 371469
rect 60625 371409 60659 371469
rect 60743 371409 60777 371469
rect 60901 371409 60935 371469
rect 61019 371409 61053 371469
rect 61177 371409 61211 371469
rect 61295 371409 61329 371469
rect 61453 371409 61487 371469
rect 61571 371409 61605 371469
rect 61729 371409 61763 371469
rect 61847 371409 61881 371469
rect 62005 371409 62039 371469
rect 62123 371409 62157 371469
rect 62281 371409 62315 371469
rect 62399 371409 62433 371469
rect 62557 371409 62591 371469
rect 62675 371409 62709 371469
rect 62833 371409 62867 371469
rect 62951 371409 62985 371469
rect 63109 371409 63143 371469
rect 63227 371409 63261 371469
rect 63385 371409 63419 371469
rect 63503 371409 63537 371469
rect 63661 371409 63695 371469
rect 63779 371409 63813 371469
rect 63937 371409 63971 371469
rect 64055 371409 64089 371469
rect 64213 371409 64247 371469
rect 64331 371409 64365 371469
rect 64489 371409 64523 371469
rect 64607 371409 64641 371469
rect 64765 371409 64799 371469
rect 64883 371409 64917 371469
rect 65041 371409 65075 371469
rect 65159 371409 65193 371469
rect 65317 371409 65351 371469
rect 65435 371409 65469 371469
rect 65593 371409 65627 371469
rect 65711 371409 65745 371469
rect 65869 371409 65903 371469
rect 65987 371409 66021 371469
rect 66145 371409 66179 371469
rect 66263 371409 66297 371469
rect 66421 371409 66455 371469
rect 66539 371409 66573 371469
rect 66697 371409 66731 371469
rect 66815 371409 66849 371469
rect 66973 371409 67007 371469
rect 67091 371409 67125 371469
rect 67249 371409 67283 371469
rect 53353 371325 53421 371359
rect 53629 371325 53697 371359
rect 53905 371325 53973 371359
rect 54181 371325 54249 371359
rect 54457 371325 54525 371359
rect 54733 371325 54801 371359
rect 55009 371325 55077 371359
rect 55285 371325 55353 371359
rect 55561 371325 55629 371359
rect 55837 371325 55905 371359
rect 56113 371325 56181 371359
rect 56389 371325 56457 371359
rect 56665 371325 56733 371359
rect 56941 371325 57009 371359
rect 57217 371325 57285 371359
rect 57493 371325 57561 371359
rect 57769 371325 57837 371359
rect 58045 371325 58113 371359
rect 58321 371325 58389 371359
rect 58597 371325 58665 371359
rect 58873 371325 58941 371359
rect 59149 371325 59217 371359
rect 59425 371325 59493 371359
rect 59701 371325 59769 371359
rect 59977 371325 60045 371359
rect 60253 371325 60321 371359
rect 60529 371325 60597 371359
rect 60805 371325 60873 371359
rect 61081 371325 61149 371359
rect 61357 371325 61425 371359
rect 61633 371325 61701 371359
rect 61909 371325 61977 371359
rect 62185 371325 62253 371359
rect 62461 371325 62529 371359
rect 62737 371325 62805 371359
rect 63013 371325 63081 371359
rect 63289 371325 63357 371359
rect 63565 371325 63633 371359
rect 63841 371325 63909 371359
rect 64117 371325 64185 371359
rect 64393 371325 64461 371359
rect 64669 371325 64737 371359
rect 64945 371325 65013 371359
rect 65221 371325 65289 371359
rect 65497 371325 65565 371359
rect 65773 371325 65841 371359
rect 66049 371325 66117 371359
rect 66325 371325 66393 371359
rect 66601 371325 66669 371359
rect 66877 371325 66945 371359
rect 67153 371325 67221 371359
rect 143353 371519 143421 371553
rect 143629 371519 143697 371553
rect 143905 371519 143973 371553
rect 144181 371519 144249 371553
rect 144457 371519 144525 371553
rect 144733 371519 144801 371553
rect 145009 371519 145077 371553
rect 145285 371519 145353 371553
rect 145561 371519 145629 371553
rect 145837 371519 145905 371553
rect 146113 371519 146181 371553
rect 146389 371519 146457 371553
rect 146665 371519 146733 371553
rect 146941 371519 147009 371553
rect 147217 371519 147285 371553
rect 147493 371519 147561 371553
rect 147769 371519 147837 371553
rect 148045 371519 148113 371553
rect 148321 371519 148389 371553
rect 148597 371519 148665 371553
rect 148873 371519 148941 371553
rect 149149 371519 149217 371553
rect 149425 371519 149493 371553
rect 149701 371519 149769 371553
rect 149977 371519 150045 371553
rect 150253 371519 150321 371553
rect 150529 371519 150597 371553
rect 150805 371519 150873 371553
rect 151081 371519 151149 371553
rect 151357 371519 151425 371553
rect 151633 371519 151701 371553
rect 151909 371519 151977 371553
rect 152185 371519 152253 371553
rect 152461 371519 152529 371553
rect 152737 371519 152805 371553
rect 153013 371519 153081 371553
rect 153289 371519 153357 371553
rect 153565 371519 153633 371553
rect 153841 371519 153909 371553
rect 154117 371519 154185 371553
rect 154393 371519 154461 371553
rect 154669 371519 154737 371553
rect 154945 371519 155013 371553
rect 155221 371519 155289 371553
rect 155497 371519 155565 371553
rect 155773 371519 155841 371553
rect 156049 371519 156117 371553
rect 156325 371519 156393 371553
rect 156601 371519 156669 371553
rect 156877 371519 156945 371553
rect 157153 371519 157221 371553
rect 143291 371409 143325 371469
rect 143449 371409 143483 371469
rect 143567 371409 143601 371469
rect 143725 371409 143759 371469
rect 143843 371409 143877 371469
rect 144001 371409 144035 371469
rect 144119 371409 144153 371469
rect 144277 371409 144311 371469
rect 144395 371409 144429 371469
rect 144553 371409 144587 371469
rect 144671 371409 144705 371469
rect 144829 371409 144863 371469
rect 144947 371409 144981 371469
rect 145105 371409 145139 371469
rect 145223 371409 145257 371469
rect 145381 371409 145415 371469
rect 145499 371409 145533 371469
rect 145657 371409 145691 371469
rect 145775 371409 145809 371469
rect 145933 371409 145967 371469
rect 146051 371409 146085 371469
rect 146209 371409 146243 371469
rect 146327 371409 146361 371469
rect 146485 371409 146519 371469
rect 146603 371409 146637 371469
rect 146761 371409 146795 371469
rect 146879 371409 146913 371469
rect 147037 371409 147071 371469
rect 147155 371409 147189 371469
rect 147313 371409 147347 371469
rect 147431 371409 147465 371469
rect 147589 371409 147623 371469
rect 147707 371409 147741 371469
rect 147865 371409 147899 371469
rect 147983 371409 148017 371469
rect 148141 371409 148175 371469
rect 148259 371409 148293 371469
rect 148417 371409 148451 371469
rect 148535 371409 148569 371469
rect 148693 371409 148727 371469
rect 148811 371409 148845 371469
rect 148969 371409 149003 371469
rect 149087 371409 149121 371469
rect 149245 371409 149279 371469
rect 149363 371409 149397 371469
rect 149521 371409 149555 371469
rect 149639 371409 149673 371469
rect 149797 371409 149831 371469
rect 149915 371409 149949 371469
rect 150073 371409 150107 371469
rect 150191 371409 150225 371469
rect 150349 371409 150383 371469
rect 150467 371409 150501 371469
rect 150625 371409 150659 371469
rect 150743 371409 150777 371469
rect 150901 371409 150935 371469
rect 151019 371409 151053 371469
rect 151177 371409 151211 371469
rect 151295 371409 151329 371469
rect 151453 371409 151487 371469
rect 151571 371409 151605 371469
rect 151729 371409 151763 371469
rect 151847 371409 151881 371469
rect 152005 371409 152039 371469
rect 152123 371409 152157 371469
rect 152281 371409 152315 371469
rect 152399 371409 152433 371469
rect 152557 371409 152591 371469
rect 152675 371409 152709 371469
rect 152833 371409 152867 371469
rect 152951 371409 152985 371469
rect 153109 371409 153143 371469
rect 153227 371409 153261 371469
rect 153385 371409 153419 371469
rect 153503 371409 153537 371469
rect 153661 371409 153695 371469
rect 153779 371409 153813 371469
rect 153937 371409 153971 371469
rect 154055 371409 154089 371469
rect 154213 371409 154247 371469
rect 154331 371409 154365 371469
rect 154489 371409 154523 371469
rect 154607 371409 154641 371469
rect 154765 371409 154799 371469
rect 154883 371409 154917 371469
rect 155041 371409 155075 371469
rect 155159 371409 155193 371469
rect 155317 371409 155351 371469
rect 155435 371409 155469 371469
rect 155593 371409 155627 371469
rect 155711 371409 155745 371469
rect 155869 371409 155903 371469
rect 155987 371409 156021 371469
rect 156145 371409 156179 371469
rect 156263 371409 156297 371469
rect 156421 371409 156455 371469
rect 156539 371409 156573 371469
rect 156697 371409 156731 371469
rect 156815 371409 156849 371469
rect 156973 371409 157007 371469
rect 157091 371409 157125 371469
rect 157249 371409 157283 371469
rect 143353 371325 143421 371359
rect 143629 371325 143697 371359
rect 143905 371325 143973 371359
rect 144181 371325 144249 371359
rect 144457 371325 144525 371359
rect 144733 371325 144801 371359
rect 145009 371325 145077 371359
rect 145285 371325 145353 371359
rect 145561 371325 145629 371359
rect 145837 371325 145905 371359
rect 146113 371325 146181 371359
rect 146389 371325 146457 371359
rect 146665 371325 146733 371359
rect 146941 371325 147009 371359
rect 147217 371325 147285 371359
rect 147493 371325 147561 371359
rect 147769 371325 147837 371359
rect 148045 371325 148113 371359
rect 148321 371325 148389 371359
rect 148597 371325 148665 371359
rect 148873 371325 148941 371359
rect 149149 371325 149217 371359
rect 149425 371325 149493 371359
rect 149701 371325 149769 371359
rect 149977 371325 150045 371359
rect 150253 371325 150321 371359
rect 150529 371325 150597 371359
rect 150805 371325 150873 371359
rect 151081 371325 151149 371359
rect 151357 371325 151425 371359
rect 151633 371325 151701 371359
rect 151909 371325 151977 371359
rect 152185 371325 152253 371359
rect 152461 371325 152529 371359
rect 152737 371325 152805 371359
rect 153013 371325 153081 371359
rect 153289 371325 153357 371359
rect 153565 371325 153633 371359
rect 153841 371325 153909 371359
rect 154117 371325 154185 371359
rect 154393 371325 154461 371359
rect 154669 371325 154737 371359
rect 154945 371325 155013 371359
rect 155221 371325 155289 371359
rect 155497 371325 155565 371359
rect 155773 371325 155841 371359
rect 156049 371325 156117 371359
rect 156325 371325 156393 371359
rect 156601 371325 156669 371359
rect 156877 371325 156945 371359
rect 157153 371325 157221 371359
rect 334933 372003 335001 372037
rect 335209 372003 335277 372037
rect 335485 372003 335553 372037
rect 335761 372003 335829 372037
rect 336037 372003 336105 372037
rect 336313 372003 336381 372037
rect 336589 372003 336657 372037
rect 336865 372003 336933 372037
rect 337141 372003 337209 372037
rect 337417 372003 337485 372037
rect 337693 372003 337761 372037
rect 327886 371706 327964 371762
rect 323904 371644 323958 371686
rect 418903 371809 418971 371843
rect 419179 371809 419247 371843
rect 419455 371809 419523 371843
rect 419731 371809 419799 371843
rect 420007 371809 420075 371843
rect 420283 371809 420351 371843
rect 420559 371809 420627 371843
rect 420835 371809 420903 371843
rect 421111 371809 421179 371843
rect 421387 371809 421455 371843
rect 418841 371699 418875 371759
rect 418999 371699 419033 371759
rect 419117 371699 419151 371759
rect 419275 371699 419309 371759
rect 419393 371699 419427 371759
rect 419551 371699 419585 371759
rect 419669 371699 419703 371759
rect 419827 371699 419861 371759
rect 419945 371699 419979 371759
rect 420103 371699 420137 371759
rect 420221 371699 420255 371759
rect 420379 371699 420413 371759
rect 420497 371699 420531 371759
rect 420655 371699 420689 371759
rect 420773 371699 420807 371759
rect 420931 371699 420965 371759
rect 421049 371699 421083 371759
rect 421207 371699 421241 371759
rect 421325 371699 421359 371759
rect 421483 371699 421517 371759
rect 418903 371615 418971 371649
rect 419179 371615 419247 371649
rect 419455 371615 419523 371649
rect 419731 371615 419799 371649
rect 420007 371615 420075 371649
rect 420283 371615 420351 371649
rect 420559 371615 420627 371649
rect 420835 371615 420903 371649
rect 421111 371615 421179 371649
rect 421387 371615 421455 371649
rect 419566 371290 419638 371334
rect 508902 371481 508970 371515
rect 509178 371481 509246 371515
rect 509454 371481 509522 371515
rect 509730 371481 509798 371515
rect 510006 371481 510074 371515
rect 508840 371371 508874 371431
rect 508998 371371 509032 371431
rect 509116 371371 509150 371431
rect 509274 371371 509308 371431
rect 509392 371371 509426 371431
rect 509550 371371 509584 371431
rect 509668 371371 509702 371431
rect 509826 371371 509860 371431
rect 509944 371371 509978 371431
rect 510102 371371 510136 371431
rect 508902 371287 508970 371321
rect 509178 371287 509246 371321
rect 509454 371287 509522 371321
rect 509730 371287 509798 371321
rect 510006 371287 510074 371321
rect 508923 371210 508961 371244
rect 57346 371029 57424 371085
rect 147346 371029 147424 371085
rect 232710 370923 232778 370957
rect 232986 370923 233054 370957
rect 233262 370923 233330 370957
rect 233538 370923 233606 370957
rect 233814 370923 233882 370957
rect 234090 370923 234158 370957
rect 234366 370923 234434 370957
rect 234642 370923 234710 370957
rect 234918 370923 234986 370957
rect 235194 370923 235262 370957
rect 235470 370923 235538 370957
rect 235746 370923 235814 370957
rect 236022 370923 236090 370957
rect 236298 370923 236366 370957
rect 236574 370923 236642 370957
rect 236850 370923 236918 370957
rect 237126 370923 237194 370957
rect 237402 370923 237470 370957
rect 237678 370923 237746 370957
rect 237954 370923 238022 370957
rect 238230 370923 238298 370957
rect 238506 370923 238574 370957
rect 238782 370923 238850 370957
rect 239058 370923 239126 370957
rect 239334 370923 239402 370957
rect 239610 370923 239678 370957
rect 239886 370923 239954 370957
rect 240162 370923 240230 370957
rect 240438 370923 240506 370957
rect 240714 370923 240782 370957
rect 240990 370923 241058 370957
rect 241266 370923 241334 370957
rect 241542 370923 241610 370957
rect 241818 370923 241886 370957
rect 242094 370923 242162 370957
rect 242370 370923 242438 370957
rect 242646 370923 242714 370957
rect 242922 370923 242990 370957
rect 243198 370923 243266 370957
rect 243474 370923 243542 370957
rect 243750 370923 243818 370957
rect 244026 370923 244094 370957
rect 244302 370923 244370 370957
rect 244578 370923 244646 370957
rect 244854 370923 244922 370957
rect 245130 370923 245198 370957
rect 245406 370923 245474 370957
rect 245682 370923 245750 370957
rect 245958 370923 246026 370957
rect 246234 370923 246302 370957
rect 246510 370923 246578 370957
rect 232648 370813 232682 370873
rect 232806 370813 232840 370873
rect 232924 370813 232958 370873
rect 233082 370813 233116 370873
rect 233200 370813 233234 370873
rect 233358 370813 233392 370873
rect 233476 370813 233510 370873
rect 233634 370813 233668 370873
rect 233752 370813 233786 370873
rect 233910 370813 233944 370873
rect 234028 370813 234062 370873
rect 234186 370813 234220 370873
rect 234304 370813 234338 370873
rect 234462 370813 234496 370873
rect 234580 370813 234614 370873
rect 234738 370813 234772 370873
rect 234856 370813 234890 370873
rect 235014 370813 235048 370873
rect 235132 370813 235166 370873
rect 235290 370813 235324 370873
rect 235408 370813 235442 370873
rect 235566 370813 235600 370873
rect 235684 370813 235718 370873
rect 235842 370813 235876 370873
rect 235960 370813 235994 370873
rect 236118 370813 236152 370873
rect 236236 370813 236270 370873
rect 236394 370813 236428 370873
rect 236512 370813 236546 370873
rect 236670 370813 236704 370873
rect 236788 370813 236822 370873
rect 236946 370813 236980 370873
rect 237064 370813 237098 370873
rect 237222 370813 237256 370873
rect 237340 370813 237374 370873
rect 237498 370813 237532 370873
rect 237616 370813 237650 370873
rect 237774 370813 237808 370873
rect 237892 370813 237926 370873
rect 238050 370813 238084 370873
rect 238168 370813 238202 370873
rect 238326 370813 238360 370873
rect 238444 370813 238478 370873
rect 238602 370813 238636 370873
rect 238720 370813 238754 370873
rect 238878 370813 238912 370873
rect 238996 370813 239030 370873
rect 239154 370813 239188 370873
rect 239272 370813 239306 370873
rect 239430 370813 239464 370873
rect 239548 370813 239582 370873
rect 239706 370813 239740 370873
rect 239824 370813 239858 370873
rect 239982 370813 240016 370873
rect 240100 370813 240134 370873
rect 240258 370813 240292 370873
rect 240376 370813 240410 370873
rect 240534 370813 240568 370873
rect 240652 370813 240686 370873
rect 240810 370813 240844 370873
rect 240928 370813 240962 370873
rect 241086 370813 241120 370873
rect 241204 370813 241238 370873
rect 241362 370813 241396 370873
rect 241480 370813 241514 370873
rect 241638 370813 241672 370873
rect 241756 370813 241790 370873
rect 241914 370813 241948 370873
rect 242032 370813 242066 370873
rect 242190 370813 242224 370873
rect 242308 370813 242342 370873
rect 242466 370813 242500 370873
rect 242584 370813 242618 370873
rect 242742 370813 242776 370873
rect 242860 370813 242894 370873
rect 243018 370813 243052 370873
rect 243136 370813 243170 370873
rect 243294 370813 243328 370873
rect 243412 370813 243446 370873
rect 243570 370813 243604 370873
rect 243688 370813 243722 370873
rect 243846 370813 243880 370873
rect 243964 370813 243998 370873
rect 244122 370813 244156 370873
rect 244240 370813 244274 370873
rect 244398 370813 244432 370873
rect 244516 370813 244550 370873
rect 244674 370813 244708 370873
rect 244792 370813 244826 370873
rect 244950 370813 244984 370873
rect 245068 370813 245102 370873
rect 245226 370813 245260 370873
rect 245344 370813 245378 370873
rect 245502 370813 245536 370873
rect 245620 370813 245654 370873
rect 245778 370813 245812 370873
rect 245896 370813 245930 370873
rect 246054 370813 246088 370873
rect 246172 370813 246206 370873
rect 246330 370813 246364 370873
rect 246448 370813 246482 370873
rect 246606 370813 246640 370873
rect 232710 370729 232778 370763
rect 232986 370729 233054 370763
rect 233262 370729 233330 370763
rect 233538 370729 233606 370763
rect 233814 370729 233882 370763
rect 234090 370729 234158 370763
rect 234366 370729 234434 370763
rect 234642 370729 234710 370763
rect 234918 370729 234986 370763
rect 235194 370729 235262 370763
rect 235470 370729 235538 370763
rect 235746 370729 235814 370763
rect 236022 370729 236090 370763
rect 236298 370729 236366 370763
rect 236574 370729 236642 370763
rect 236850 370729 236918 370763
rect 237126 370729 237194 370763
rect 237402 370729 237470 370763
rect 237678 370729 237746 370763
rect 237954 370729 238022 370763
rect 238230 370729 238298 370763
rect 238506 370729 238574 370763
rect 238782 370729 238850 370763
rect 239058 370729 239126 370763
rect 239334 370729 239402 370763
rect 239610 370729 239678 370763
rect 239886 370729 239954 370763
rect 240162 370729 240230 370763
rect 240438 370729 240506 370763
rect 240714 370729 240782 370763
rect 240990 370729 241058 370763
rect 241266 370729 241334 370763
rect 241542 370729 241610 370763
rect 241818 370729 241886 370763
rect 242094 370729 242162 370763
rect 242370 370729 242438 370763
rect 242646 370729 242714 370763
rect 242922 370729 242990 370763
rect 243198 370729 243266 370763
rect 243474 370729 243542 370763
rect 243750 370729 243818 370763
rect 244026 370729 244094 370763
rect 244302 370729 244370 370763
rect 244578 370729 244646 370763
rect 244854 370729 244922 370763
rect 245130 370729 245198 370763
rect 245406 370729 245474 370763
rect 245682 370729 245750 370763
rect 245958 370729 246026 370763
rect 246234 370729 246302 370763
rect 246510 370729 246578 370763
rect 236703 370433 236781 370489
rect 234282 252164 234336 252206
rect 234271 251805 234339 251839
rect 234547 251805 234615 251839
rect 234823 251805 234891 251839
rect 235099 251805 235167 251839
rect 235375 251805 235443 251839
rect 235651 251805 235719 251839
rect 235927 251805 235995 251839
rect 236203 251805 236271 251839
rect 236479 251805 236547 251839
rect 236755 251805 236823 251839
rect 237031 251805 237099 251839
rect 237307 251805 237375 251839
rect 237583 251805 237651 251839
rect 237859 251805 237927 251839
rect 238135 251805 238203 251839
rect 238411 251805 238479 251839
rect 238687 251805 238755 251839
rect 238963 251805 239031 251839
rect 239239 251805 239307 251839
rect 239515 251805 239583 251839
rect 239791 251805 239859 251839
rect 240067 251805 240135 251839
rect 240343 251805 240411 251839
rect 240619 251805 240687 251839
rect 240895 251805 240963 251839
rect 241171 251805 241239 251839
rect 241447 251805 241515 251839
rect 241723 251805 241791 251839
rect 241999 251805 242067 251839
rect 242275 251805 242343 251839
rect 242551 251805 242619 251839
rect 242827 251805 242895 251839
rect 243103 251805 243171 251839
rect 243379 251805 243447 251839
rect 243655 251805 243723 251839
rect 243931 251805 243999 251839
rect 244207 251805 244275 251839
rect 244483 251805 244551 251839
rect 244759 251805 244827 251839
rect 245035 251805 245103 251839
rect 245311 251805 245379 251839
rect 245587 251805 245655 251839
rect 245863 251805 245931 251839
rect 246139 251805 246207 251839
rect 246415 251805 246483 251839
rect 246691 251805 246759 251839
rect 246967 251805 247035 251839
rect 247243 251805 247311 251839
rect 247519 251805 247587 251839
rect 247795 251805 247863 251839
rect 248071 251805 248139 251839
rect 58902 251481 58970 251515
rect 59178 251481 59246 251515
rect 59454 251481 59522 251515
rect 59730 251481 59798 251515
rect 60006 251481 60074 251515
rect 58840 251371 58874 251431
rect 58998 251371 59032 251431
rect 59116 251371 59150 251431
rect 59274 251371 59308 251431
rect 59392 251371 59426 251431
rect 59550 251371 59584 251431
rect 59668 251371 59702 251431
rect 59826 251371 59860 251431
rect 59944 251371 59978 251431
rect 60102 251371 60136 251431
rect 58902 251287 58970 251321
rect 59178 251287 59246 251321
rect 59454 251287 59522 251321
rect 59730 251287 59798 251321
rect 60006 251287 60074 251321
rect 58923 251210 58961 251244
rect 148027 251605 148095 251639
rect 148303 251605 148371 251639
rect 148579 251605 148647 251639
rect 148855 251605 148923 251639
rect 149131 251605 149199 251639
rect 149407 251605 149475 251639
rect 149683 251605 149751 251639
rect 149959 251605 150027 251639
rect 150235 251605 150303 251639
rect 150511 251605 150579 251639
rect 147965 251495 147999 251555
rect 148123 251495 148157 251555
rect 148241 251495 148275 251555
rect 148399 251495 148433 251555
rect 148517 251495 148551 251555
rect 148675 251495 148709 251555
rect 148793 251495 148827 251555
rect 148951 251495 148985 251555
rect 149069 251495 149103 251555
rect 149227 251495 149261 251555
rect 149345 251495 149379 251555
rect 149503 251495 149537 251555
rect 149621 251495 149655 251555
rect 149779 251495 149813 251555
rect 149897 251495 149931 251555
rect 150055 251495 150089 251555
rect 150173 251495 150207 251555
rect 150331 251495 150365 251555
rect 150449 251495 150483 251555
rect 150607 251495 150641 251555
rect 148027 251411 148095 251445
rect 148303 251411 148371 251445
rect 148579 251411 148647 251445
rect 148855 251411 148923 251445
rect 149131 251411 149199 251445
rect 149407 251411 149475 251445
rect 149683 251411 149751 251445
rect 149959 251411 150027 251445
rect 150235 251411 150303 251445
rect 150511 251411 150579 251445
rect 234209 251695 234243 251755
rect 234367 251695 234401 251755
rect 234485 251695 234519 251755
rect 234643 251695 234677 251755
rect 234761 251695 234795 251755
rect 234919 251695 234953 251755
rect 235037 251695 235071 251755
rect 235195 251695 235229 251755
rect 235313 251695 235347 251755
rect 235471 251695 235505 251755
rect 235589 251695 235623 251755
rect 235747 251695 235781 251755
rect 235865 251695 235899 251755
rect 236023 251695 236057 251755
rect 236141 251695 236175 251755
rect 236299 251695 236333 251755
rect 236417 251695 236451 251755
rect 236575 251695 236609 251755
rect 236693 251695 236727 251755
rect 236851 251695 236885 251755
rect 236969 251695 237003 251755
rect 237127 251695 237161 251755
rect 237245 251695 237279 251755
rect 237403 251695 237437 251755
rect 237521 251695 237555 251755
rect 237679 251695 237713 251755
rect 237797 251695 237831 251755
rect 237955 251695 237989 251755
rect 238073 251695 238107 251755
rect 238231 251695 238265 251755
rect 238349 251695 238383 251755
rect 238507 251695 238541 251755
rect 238625 251695 238659 251755
rect 238783 251695 238817 251755
rect 238901 251695 238935 251755
rect 239059 251695 239093 251755
rect 239177 251695 239211 251755
rect 239335 251695 239369 251755
rect 239453 251695 239487 251755
rect 239611 251695 239645 251755
rect 239729 251695 239763 251755
rect 239887 251695 239921 251755
rect 240005 251695 240039 251755
rect 240163 251695 240197 251755
rect 240281 251695 240315 251755
rect 240439 251695 240473 251755
rect 240557 251695 240591 251755
rect 240715 251695 240749 251755
rect 240833 251695 240867 251755
rect 240991 251695 241025 251755
rect 241109 251695 241143 251755
rect 241267 251695 241301 251755
rect 241385 251695 241419 251755
rect 241543 251695 241577 251755
rect 241661 251695 241695 251755
rect 241819 251695 241853 251755
rect 241937 251695 241971 251755
rect 242095 251695 242129 251755
rect 242213 251695 242247 251755
rect 242371 251695 242405 251755
rect 242489 251695 242523 251755
rect 242647 251695 242681 251755
rect 242765 251695 242799 251755
rect 242923 251695 242957 251755
rect 243041 251695 243075 251755
rect 243199 251695 243233 251755
rect 243317 251695 243351 251755
rect 243475 251695 243509 251755
rect 243593 251695 243627 251755
rect 243751 251695 243785 251755
rect 243869 251695 243903 251755
rect 244027 251695 244061 251755
rect 244145 251695 244179 251755
rect 244303 251695 244337 251755
rect 244421 251695 244455 251755
rect 244579 251695 244613 251755
rect 244697 251695 244731 251755
rect 244855 251695 244889 251755
rect 244973 251695 245007 251755
rect 245131 251695 245165 251755
rect 245249 251695 245283 251755
rect 245407 251695 245441 251755
rect 245525 251695 245559 251755
rect 245683 251695 245717 251755
rect 245801 251695 245835 251755
rect 245959 251695 245993 251755
rect 246077 251695 246111 251755
rect 246235 251695 246269 251755
rect 246353 251695 246387 251755
rect 246511 251695 246545 251755
rect 246629 251695 246663 251755
rect 246787 251695 246821 251755
rect 246905 251695 246939 251755
rect 247063 251695 247097 251755
rect 247181 251695 247215 251755
rect 247339 251695 247373 251755
rect 247457 251695 247491 251755
rect 247615 251695 247649 251755
rect 247733 251695 247767 251755
rect 247891 251695 247925 251755
rect 248009 251695 248043 251755
rect 248167 251695 248201 251755
rect 234271 251611 234339 251645
rect 234547 251611 234615 251645
rect 234823 251611 234891 251645
rect 235099 251611 235167 251645
rect 235375 251611 235443 251645
rect 235651 251611 235719 251645
rect 235927 251611 235995 251645
rect 236203 251611 236271 251645
rect 236479 251611 236547 251645
rect 236755 251611 236823 251645
rect 237031 251611 237099 251645
rect 237307 251611 237375 251645
rect 237583 251611 237651 251645
rect 237859 251611 237927 251645
rect 238135 251611 238203 251645
rect 238411 251611 238479 251645
rect 238687 251611 238755 251645
rect 238963 251611 239031 251645
rect 239239 251611 239307 251645
rect 239515 251611 239583 251645
rect 239791 251611 239859 251645
rect 240067 251611 240135 251645
rect 240343 251611 240411 251645
rect 240619 251611 240687 251645
rect 240895 251611 240963 251645
rect 241171 251611 241239 251645
rect 241447 251611 241515 251645
rect 241723 251611 241791 251645
rect 241999 251611 242067 251645
rect 242275 251611 242343 251645
rect 242551 251611 242619 251645
rect 242827 251611 242895 251645
rect 243103 251611 243171 251645
rect 243379 251611 243447 251645
rect 243655 251611 243723 251645
rect 243931 251611 243999 251645
rect 244207 251611 244275 251645
rect 244483 251611 244551 251645
rect 244759 251611 244827 251645
rect 245035 251611 245103 251645
rect 245311 251611 245379 251645
rect 245587 251611 245655 251645
rect 245863 251611 245931 251645
rect 246139 251611 246207 251645
rect 246415 251611 246483 251645
rect 246691 251611 246759 251645
rect 246967 251611 247035 251645
rect 247243 251611 247311 251645
rect 247519 251611 247587 251645
rect 247795 251611 247863 251645
rect 248071 251611 248139 251645
rect 413353 251519 413421 251553
rect 413629 251519 413697 251553
rect 413905 251519 413973 251553
rect 414181 251519 414249 251553
rect 414457 251519 414525 251553
rect 414733 251519 414801 251553
rect 415009 251519 415077 251553
rect 415285 251519 415353 251553
rect 415561 251519 415629 251553
rect 415837 251519 415905 251553
rect 416113 251519 416181 251553
rect 416389 251519 416457 251553
rect 416665 251519 416733 251553
rect 416941 251519 417009 251553
rect 417217 251519 417285 251553
rect 417493 251519 417561 251553
rect 417769 251519 417837 251553
rect 418045 251519 418113 251553
rect 418321 251519 418389 251553
rect 418597 251519 418665 251553
rect 418873 251519 418941 251553
rect 419149 251519 419217 251553
rect 419425 251519 419493 251553
rect 419701 251519 419769 251553
rect 419977 251519 420045 251553
rect 420253 251519 420321 251553
rect 420529 251519 420597 251553
rect 420805 251519 420873 251553
rect 421081 251519 421149 251553
rect 421357 251519 421425 251553
rect 421633 251519 421701 251553
rect 421909 251519 421977 251553
rect 422185 251519 422253 251553
rect 422461 251519 422529 251553
rect 422737 251519 422805 251553
rect 423013 251519 423081 251553
rect 423289 251519 423357 251553
rect 423565 251519 423633 251553
rect 423841 251519 423909 251553
rect 424117 251519 424185 251553
rect 424393 251519 424461 251553
rect 424669 251519 424737 251553
rect 424945 251519 425013 251553
rect 425221 251519 425289 251553
rect 425497 251519 425565 251553
rect 425773 251519 425841 251553
rect 426049 251519 426117 251553
rect 426325 251519 426393 251553
rect 426601 251519 426669 251553
rect 426877 251519 426945 251553
rect 427153 251519 427221 251553
rect 413291 251409 413325 251469
rect 413449 251409 413483 251469
rect 413567 251409 413601 251469
rect 413725 251409 413759 251469
rect 413843 251409 413877 251469
rect 414001 251409 414035 251469
rect 414119 251409 414153 251469
rect 414277 251409 414311 251469
rect 414395 251409 414429 251469
rect 414553 251409 414587 251469
rect 414671 251409 414705 251469
rect 414829 251409 414863 251469
rect 414947 251409 414981 251469
rect 415105 251409 415139 251469
rect 415223 251409 415257 251469
rect 415381 251409 415415 251469
rect 415499 251409 415533 251469
rect 415657 251409 415691 251469
rect 415775 251409 415809 251469
rect 415933 251409 415967 251469
rect 416051 251409 416085 251469
rect 416209 251409 416243 251469
rect 416327 251409 416361 251469
rect 416485 251409 416519 251469
rect 416603 251409 416637 251469
rect 416761 251409 416795 251469
rect 416879 251409 416913 251469
rect 417037 251409 417071 251469
rect 417155 251409 417189 251469
rect 417313 251409 417347 251469
rect 417431 251409 417465 251469
rect 417589 251409 417623 251469
rect 417707 251409 417741 251469
rect 417865 251409 417899 251469
rect 417983 251409 418017 251469
rect 418141 251409 418175 251469
rect 418259 251409 418293 251469
rect 418417 251409 418451 251469
rect 418535 251409 418569 251469
rect 418693 251409 418727 251469
rect 418811 251409 418845 251469
rect 418969 251409 419003 251469
rect 419087 251409 419121 251469
rect 419245 251409 419279 251469
rect 419363 251409 419397 251469
rect 419521 251409 419555 251469
rect 419639 251409 419673 251469
rect 419797 251409 419831 251469
rect 419915 251409 419949 251469
rect 420073 251409 420107 251469
rect 420191 251409 420225 251469
rect 420349 251409 420383 251469
rect 420467 251409 420501 251469
rect 420625 251409 420659 251469
rect 420743 251409 420777 251469
rect 420901 251409 420935 251469
rect 421019 251409 421053 251469
rect 421177 251409 421211 251469
rect 421295 251409 421329 251469
rect 421453 251409 421487 251469
rect 421571 251409 421605 251469
rect 421729 251409 421763 251469
rect 421847 251409 421881 251469
rect 422005 251409 422039 251469
rect 422123 251409 422157 251469
rect 422281 251409 422315 251469
rect 422399 251409 422433 251469
rect 422557 251409 422591 251469
rect 422675 251409 422709 251469
rect 422833 251409 422867 251469
rect 422951 251409 422985 251469
rect 423109 251409 423143 251469
rect 423227 251409 423261 251469
rect 423385 251409 423419 251469
rect 423503 251409 423537 251469
rect 423661 251409 423695 251469
rect 423779 251409 423813 251469
rect 423937 251409 423971 251469
rect 424055 251409 424089 251469
rect 424213 251409 424247 251469
rect 424331 251409 424365 251469
rect 424489 251409 424523 251469
rect 424607 251409 424641 251469
rect 424765 251409 424799 251469
rect 424883 251409 424917 251469
rect 425041 251409 425075 251469
rect 425159 251409 425193 251469
rect 425317 251409 425351 251469
rect 425435 251409 425469 251469
rect 425593 251409 425627 251469
rect 425711 251409 425745 251469
rect 425869 251409 425903 251469
rect 425987 251409 426021 251469
rect 426145 251409 426179 251469
rect 426263 251409 426297 251469
rect 426421 251409 426455 251469
rect 426539 251409 426573 251469
rect 426697 251409 426731 251469
rect 426815 251409 426849 251469
rect 426973 251409 427007 251469
rect 427091 251409 427125 251469
rect 427249 251409 427283 251469
rect 238264 251314 238342 251370
rect 413353 251325 413421 251359
rect 413629 251325 413697 251359
rect 413905 251325 413973 251359
rect 414181 251325 414249 251359
rect 414457 251325 414525 251359
rect 414733 251325 414801 251359
rect 415009 251325 415077 251359
rect 415285 251325 415353 251359
rect 415561 251325 415629 251359
rect 415837 251325 415905 251359
rect 416113 251325 416181 251359
rect 416389 251325 416457 251359
rect 416665 251325 416733 251359
rect 416941 251325 417009 251359
rect 417217 251325 417285 251359
rect 417493 251325 417561 251359
rect 417769 251325 417837 251359
rect 418045 251325 418113 251359
rect 418321 251325 418389 251359
rect 418597 251325 418665 251359
rect 418873 251325 418941 251359
rect 419149 251325 419217 251359
rect 419425 251325 419493 251359
rect 419701 251325 419769 251359
rect 419977 251325 420045 251359
rect 420253 251325 420321 251359
rect 420529 251325 420597 251359
rect 420805 251325 420873 251359
rect 421081 251325 421149 251359
rect 421357 251325 421425 251359
rect 421633 251325 421701 251359
rect 421909 251325 421977 251359
rect 422185 251325 422253 251359
rect 422461 251325 422529 251359
rect 422737 251325 422805 251359
rect 423013 251325 423081 251359
rect 423289 251325 423357 251359
rect 423565 251325 423633 251359
rect 423841 251325 423909 251359
rect 424117 251325 424185 251359
rect 234282 251252 234336 251294
rect 148690 251086 148762 251130
rect 322710 250923 322778 250957
rect 322986 250923 323054 250957
rect 323262 250923 323330 250957
rect 323538 250923 323606 250957
rect 323814 250923 323882 250957
rect 324090 250923 324158 250957
rect 324366 250923 324434 250957
rect 324642 250923 324710 250957
rect 324918 250923 324986 250957
rect 325194 250923 325262 250957
rect 325470 250923 325538 250957
rect 325746 250923 325814 250957
rect 326022 250923 326090 250957
rect 326298 250923 326366 250957
rect 326574 250923 326642 250957
rect 326850 250923 326918 250957
rect 327126 250923 327194 250957
rect 327402 250923 327470 250957
rect 327678 250923 327746 250957
rect 327954 250923 328022 250957
rect 328230 250923 328298 250957
rect 328506 250923 328574 250957
rect 328782 250923 328850 250957
rect 329058 250923 329126 250957
rect 329334 250923 329402 250957
rect 329610 250923 329678 250957
rect 329886 250923 329954 250957
rect 330162 250923 330230 250957
rect 330438 250923 330506 250957
rect 330714 250923 330782 250957
rect 330990 250923 331058 250957
rect 331266 250923 331334 250957
rect 331542 250923 331610 250957
rect 331818 250923 331886 250957
rect 332094 250923 332162 250957
rect 332370 250923 332438 250957
rect 332646 250923 332714 250957
rect 332922 250923 332990 250957
rect 333198 250923 333266 250957
rect 333474 250923 333542 250957
rect 333750 250923 333818 250957
rect 334026 250923 334094 250957
rect 334302 250923 334370 250957
rect 334578 250923 334646 250957
rect 334854 250923 334922 250957
rect 335130 250923 335198 250957
rect 335406 250923 335474 250957
rect 335682 250923 335750 250957
rect 335958 250923 336026 250957
rect 336234 250923 336302 250957
rect 336510 250923 336578 250957
rect 322648 250813 322682 250873
rect 322806 250813 322840 250873
rect 322924 250813 322958 250873
rect 323082 250813 323116 250873
rect 323200 250813 323234 250873
rect 323358 250813 323392 250873
rect 323476 250813 323510 250873
rect 323634 250813 323668 250873
rect 323752 250813 323786 250873
rect 323910 250813 323944 250873
rect 324028 250813 324062 250873
rect 324186 250813 324220 250873
rect 324304 250813 324338 250873
rect 324462 250813 324496 250873
rect 324580 250813 324614 250873
rect 324738 250813 324772 250873
rect 324856 250813 324890 250873
rect 325014 250813 325048 250873
rect 325132 250813 325166 250873
rect 325290 250813 325324 250873
rect 325408 250813 325442 250873
rect 325566 250813 325600 250873
rect 325684 250813 325718 250873
rect 325842 250813 325876 250873
rect 325960 250813 325994 250873
rect 326118 250813 326152 250873
rect 326236 250813 326270 250873
rect 326394 250813 326428 250873
rect 326512 250813 326546 250873
rect 326670 250813 326704 250873
rect 326788 250813 326822 250873
rect 326946 250813 326980 250873
rect 327064 250813 327098 250873
rect 327222 250813 327256 250873
rect 327340 250813 327374 250873
rect 327498 250813 327532 250873
rect 327616 250813 327650 250873
rect 327774 250813 327808 250873
rect 327892 250813 327926 250873
rect 328050 250813 328084 250873
rect 328168 250813 328202 250873
rect 328326 250813 328360 250873
rect 328444 250813 328478 250873
rect 328602 250813 328636 250873
rect 328720 250813 328754 250873
rect 328878 250813 328912 250873
rect 328996 250813 329030 250873
rect 329154 250813 329188 250873
rect 329272 250813 329306 250873
rect 329430 250813 329464 250873
rect 329548 250813 329582 250873
rect 329706 250813 329740 250873
rect 329824 250813 329858 250873
rect 329982 250813 330016 250873
rect 330100 250813 330134 250873
rect 330258 250813 330292 250873
rect 330376 250813 330410 250873
rect 330534 250813 330568 250873
rect 330652 250813 330686 250873
rect 330810 250813 330844 250873
rect 330928 250813 330962 250873
rect 331086 250813 331120 250873
rect 331204 250813 331238 250873
rect 331362 250813 331396 250873
rect 331480 250813 331514 250873
rect 331638 250813 331672 250873
rect 331756 250813 331790 250873
rect 331914 250813 331948 250873
rect 332032 250813 332066 250873
rect 332190 250813 332224 250873
rect 332308 250813 332342 250873
rect 332466 250813 332500 250873
rect 332584 250813 332618 250873
rect 332742 250813 332776 250873
rect 332860 250813 332894 250873
rect 333018 250813 333052 250873
rect 333136 250813 333170 250873
rect 333294 250813 333328 250873
rect 333412 250813 333446 250873
rect 333570 250813 333604 250873
rect 333688 250813 333722 250873
rect 333846 250813 333880 250873
rect 333964 250813 333998 250873
rect 334122 250813 334156 250873
rect 334240 250813 334274 250873
rect 334398 250813 334432 250873
rect 334516 250813 334550 250873
rect 334674 250813 334708 250873
rect 334792 250813 334826 250873
rect 334950 250813 334984 250873
rect 335068 250813 335102 250873
rect 335226 250813 335260 250873
rect 335344 250813 335378 250873
rect 335502 250813 335536 250873
rect 335620 250813 335654 250873
rect 335778 250813 335812 250873
rect 335896 250813 335930 250873
rect 336054 250813 336088 250873
rect 336172 250813 336206 250873
rect 336330 250813 336364 250873
rect 336448 250813 336482 250873
rect 336606 250813 336640 250873
rect 322710 250729 322778 250763
rect 322986 250729 323054 250763
rect 323262 250729 323330 250763
rect 323538 250729 323606 250763
rect 323814 250729 323882 250763
rect 324090 250729 324158 250763
rect 324366 250729 324434 250763
rect 324642 250729 324710 250763
rect 324918 250729 324986 250763
rect 325194 250729 325262 250763
rect 325470 250729 325538 250763
rect 325746 250729 325814 250763
rect 326022 250729 326090 250763
rect 326298 250729 326366 250763
rect 326574 250729 326642 250763
rect 326850 250729 326918 250763
rect 327126 250729 327194 250763
rect 327402 250729 327470 250763
rect 327678 250729 327746 250763
rect 327954 250729 328022 250763
rect 328230 250729 328298 250763
rect 328506 250729 328574 250763
rect 328782 250729 328850 250763
rect 329058 250729 329126 250763
rect 329334 250729 329402 250763
rect 329610 250729 329678 250763
rect 329886 250729 329954 250763
rect 330162 250729 330230 250763
rect 330438 250729 330506 250763
rect 330714 250729 330782 250763
rect 330990 250729 331058 250763
rect 331266 250729 331334 250763
rect 331542 250729 331610 250763
rect 331818 250729 331886 250763
rect 332094 250729 332162 250763
rect 332370 250729 332438 250763
rect 332646 250729 332714 250763
rect 332922 250729 332990 250763
rect 333198 250729 333266 250763
rect 333474 250729 333542 250763
rect 333750 250729 333818 250763
rect 334026 250729 334094 250763
rect 334302 250729 334370 250763
rect 334578 250729 334646 250763
rect 334854 250729 334922 250763
rect 335130 250729 335198 250763
rect 335406 250729 335474 250763
rect 335682 250729 335750 250763
rect 335958 250729 336026 250763
rect 336234 250729 336302 250763
rect 336510 250729 336578 250763
rect 424393 251325 424461 251359
rect 424669 251325 424737 251359
rect 424945 251325 425013 251359
rect 425221 251325 425289 251359
rect 425497 251325 425565 251359
rect 425773 251325 425841 251359
rect 426049 251325 426117 251359
rect 426325 251325 426393 251359
rect 426601 251325 426669 251359
rect 426877 251325 426945 251359
rect 427153 251325 427221 251359
rect 503353 251519 503421 251553
rect 503629 251519 503697 251553
rect 503905 251519 503973 251553
rect 504181 251519 504249 251553
rect 504457 251519 504525 251553
rect 504733 251519 504801 251553
rect 505009 251519 505077 251553
rect 505285 251519 505353 251553
rect 505561 251519 505629 251553
rect 505837 251519 505905 251553
rect 506113 251519 506181 251553
rect 506389 251519 506457 251553
rect 506665 251519 506733 251553
rect 506941 251519 507009 251553
rect 507217 251519 507285 251553
rect 507493 251519 507561 251553
rect 507769 251519 507837 251553
rect 508045 251519 508113 251553
rect 508321 251519 508389 251553
rect 508597 251519 508665 251553
rect 508873 251519 508941 251553
rect 509149 251519 509217 251553
rect 509425 251519 509493 251553
rect 509701 251519 509769 251553
rect 509977 251519 510045 251553
rect 510253 251519 510321 251553
rect 510529 251519 510597 251553
rect 510805 251519 510873 251553
rect 511081 251519 511149 251553
rect 511357 251519 511425 251553
rect 511633 251519 511701 251553
rect 511909 251519 511977 251553
rect 512185 251519 512253 251553
rect 512461 251519 512529 251553
rect 512737 251519 512805 251553
rect 513013 251519 513081 251553
rect 513289 251519 513357 251553
rect 513565 251519 513633 251553
rect 513841 251519 513909 251553
rect 514117 251519 514185 251553
rect 514393 251519 514461 251553
rect 514669 251519 514737 251553
rect 514945 251519 515013 251553
rect 515221 251519 515289 251553
rect 515497 251519 515565 251553
rect 515773 251519 515841 251553
rect 516049 251519 516117 251553
rect 516325 251519 516393 251553
rect 516601 251519 516669 251553
rect 516877 251519 516945 251553
rect 517153 251519 517221 251553
rect 503291 251409 503325 251469
rect 503449 251409 503483 251469
rect 503567 251409 503601 251469
rect 503725 251409 503759 251469
rect 503843 251409 503877 251469
rect 504001 251409 504035 251469
rect 504119 251409 504153 251469
rect 504277 251409 504311 251469
rect 504395 251409 504429 251469
rect 504553 251409 504587 251469
rect 504671 251409 504705 251469
rect 504829 251409 504863 251469
rect 504947 251409 504981 251469
rect 505105 251409 505139 251469
rect 505223 251409 505257 251469
rect 505381 251409 505415 251469
rect 505499 251409 505533 251469
rect 505657 251409 505691 251469
rect 505775 251409 505809 251469
rect 505933 251409 505967 251469
rect 506051 251409 506085 251469
rect 506209 251409 506243 251469
rect 506327 251409 506361 251469
rect 506485 251409 506519 251469
rect 506603 251409 506637 251469
rect 506761 251409 506795 251469
rect 506879 251409 506913 251469
rect 507037 251409 507071 251469
rect 507155 251409 507189 251469
rect 507313 251409 507347 251469
rect 507431 251409 507465 251469
rect 507589 251409 507623 251469
rect 507707 251409 507741 251469
rect 507865 251409 507899 251469
rect 507983 251409 508017 251469
rect 508141 251409 508175 251469
rect 508259 251409 508293 251469
rect 508417 251409 508451 251469
rect 508535 251409 508569 251469
rect 508693 251409 508727 251469
rect 508811 251409 508845 251469
rect 508969 251409 509003 251469
rect 509087 251409 509121 251469
rect 509245 251409 509279 251469
rect 509363 251409 509397 251469
rect 509521 251409 509555 251469
rect 509639 251409 509673 251469
rect 509797 251409 509831 251469
rect 509915 251409 509949 251469
rect 510073 251409 510107 251469
rect 510191 251409 510225 251469
rect 510349 251409 510383 251469
rect 510467 251409 510501 251469
rect 510625 251409 510659 251469
rect 510743 251409 510777 251469
rect 510901 251409 510935 251469
rect 511019 251409 511053 251469
rect 511177 251409 511211 251469
rect 511295 251409 511329 251469
rect 511453 251409 511487 251469
rect 511571 251409 511605 251469
rect 511729 251409 511763 251469
rect 511847 251409 511881 251469
rect 512005 251409 512039 251469
rect 512123 251409 512157 251469
rect 512281 251409 512315 251469
rect 512399 251409 512433 251469
rect 512557 251409 512591 251469
rect 512675 251409 512709 251469
rect 512833 251409 512867 251469
rect 512951 251409 512985 251469
rect 513109 251409 513143 251469
rect 513227 251409 513261 251469
rect 513385 251409 513419 251469
rect 513503 251409 513537 251469
rect 513661 251409 513695 251469
rect 513779 251409 513813 251469
rect 513937 251409 513971 251469
rect 514055 251409 514089 251469
rect 514213 251409 514247 251469
rect 514331 251409 514365 251469
rect 514489 251409 514523 251469
rect 514607 251409 514641 251469
rect 514765 251409 514799 251469
rect 514883 251409 514917 251469
rect 515041 251409 515075 251469
rect 515159 251409 515193 251469
rect 515317 251409 515351 251469
rect 515435 251409 515469 251469
rect 515593 251409 515627 251469
rect 515711 251409 515745 251469
rect 515869 251409 515903 251469
rect 515987 251409 516021 251469
rect 516145 251409 516179 251469
rect 516263 251409 516297 251469
rect 516421 251409 516455 251469
rect 516539 251409 516573 251469
rect 516697 251409 516731 251469
rect 516815 251409 516849 251469
rect 516973 251409 517007 251469
rect 517091 251409 517125 251469
rect 517249 251409 517283 251469
rect 503353 251325 503421 251359
rect 503629 251325 503697 251359
rect 503905 251325 503973 251359
rect 504181 251325 504249 251359
rect 504457 251325 504525 251359
rect 504733 251325 504801 251359
rect 505009 251325 505077 251359
rect 505285 251325 505353 251359
rect 505561 251325 505629 251359
rect 505837 251325 505905 251359
rect 506113 251325 506181 251359
rect 506389 251325 506457 251359
rect 506665 251325 506733 251359
rect 506941 251325 507009 251359
rect 507217 251325 507285 251359
rect 507493 251325 507561 251359
rect 507769 251325 507837 251359
rect 508045 251325 508113 251359
rect 508321 251325 508389 251359
rect 508597 251325 508665 251359
rect 508873 251325 508941 251359
rect 509149 251325 509217 251359
rect 509425 251325 509493 251359
rect 509701 251325 509769 251359
rect 509977 251325 510045 251359
rect 510253 251325 510321 251359
rect 510529 251325 510597 251359
rect 510805 251325 510873 251359
rect 511081 251325 511149 251359
rect 511357 251325 511425 251359
rect 511633 251325 511701 251359
rect 511909 251325 511977 251359
rect 512185 251325 512253 251359
rect 512461 251325 512529 251359
rect 512737 251325 512805 251359
rect 513013 251325 513081 251359
rect 513289 251325 513357 251359
rect 513565 251325 513633 251359
rect 513841 251325 513909 251359
rect 514117 251325 514185 251359
rect 514393 251325 514461 251359
rect 514669 251325 514737 251359
rect 514945 251325 515013 251359
rect 515221 251325 515289 251359
rect 515497 251325 515565 251359
rect 515773 251325 515841 251359
rect 516049 251325 516117 251359
rect 516325 251325 516393 251359
rect 516601 251325 516669 251359
rect 516877 251325 516945 251359
rect 517153 251325 517221 251359
rect 417346 251029 417424 251085
rect 507346 251029 507424 251085
rect 326703 250433 326781 250489
rect 59339 145993 59373 146027
rect 59295 145758 59329 145934
rect 59383 145758 59417 145934
rect 59339 145665 59373 145699
rect 239356 146022 239390 146056
rect 239312 145796 239346 145972
rect 239400 145796 239434 145972
rect 239356 145712 239390 145746
rect 329339 145993 329373 146027
rect 329295 145758 329329 145934
rect 329383 145758 329417 145934
rect 329339 145665 329373 145699
rect 149537 145589 149605 145623
rect 149475 145354 149509 145530
rect 149633 145354 149667 145530
rect 149537 145261 149605 145295
rect 509356 146022 509390 146056
rect 509312 145796 509346 145972
rect 509400 145796 509434 145972
rect 509356 145712 509390 145746
rect 419537 145589 419605 145623
rect 419475 145354 419509 145530
rect 419633 145354 419667 145530
rect 419537 145261 419605 145295
rect 59356 56022 59390 56056
rect 59312 55796 59346 55972
rect 59400 55796 59434 55972
rect 59356 55712 59390 55746
rect 149627 56021 149695 56055
rect 149565 55795 149599 55971
rect 149723 55795 149757 55971
rect 149627 55711 149695 55745
rect 329356 56022 329390 56056
rect 239637 55731 239705 55765
rect 239575 55505 239609 55681
rect 239733 55505 239767 55681
rect 239637 55421 239705 55455
rect 329312 55796 329346 55972
rect 329400 55796 329434 55972
rect 329356 55712 329390 55746
rect 419627 56021 419695 56055
rect 419565 55795 419599 55971
rect 419723 55795 419757 55971
rect 419627 55711 419695 55745
rect 509637 55731 509705 55765
rect 509575 55505 509609 55681
rect 509733 55505 509767 55681
rect 509637 55421 509705 55455
<< metal1 >>
rect 326940 661224 327900 661384
rect 326940 660624 327100 661224
rect 327700 660624 327900 661224
rect 326940 659704 327900 660624
rect 330660 661224 331620 661384
rect 330660 660624 330820 661224
rect 331420 660624 331620 661224
rect 330660 659704 331620 660624
rect 57138 659300 58098 659460
rect 57138 658700 57298 659300
rect 57898 658700 58098 659300
rect 57138 657780 58098 658700
rect 60858 659300 61818 659460
rect 60858 658700 61018 659300
rect 61618 658700 61818 659300
rect 59198 657780 59498 657790
rect 60858 657780 61818 658700
rect 57138 657190 61818 657780
rect 57138 657180 59238 657190
rect 59498 657180 61818 657190
rect 147138 659300 148098 659460
rect 147138 658700 147298 659300
rect 147898 658700 148098 659300
rect 147138 657780 148098 658700
rect 150858 659300 151818 659460
rect 150858 658700 151018 659300
rect 151618 658700 151818 659300
rect 150858 657780 151818 658700
rect 147138 657180 151818 657780
rect 237138 659300 238098 659460
rect 237138 658700 237298 659300
rect 237898 658700 238098 659300
rect 237138 657780 238098 658700
rect 240858 659300 241818 659460
rect 240858 658700 241018 659300
rect 241618 658700 241818 659300
rect 326940 659104 331620 659704
rect 416940 661224 417900 661384
rect 416940 660624 417100 661224
rect 417700 660624 417900 661224
rect 416940 659704 417900 660624
rect 420660 661224 421620 661384
rect 420660 660624 420820 661224
rect 421420 660624 421620 661224
rect 420660 659704 421620 660624
rect 416940 659104 421620 659704
rect 506940 661224 507900 661384
rect 506940 660624 507100 661224
rect 507700 660624 507900 661224
rect 506940 659704 507900 660624
rect 510660 661224 511620 661384
rect 510660 660624 510820 661224
rect 511420 660624 511620 661224
rect 510660 659704 511620 660624
rect 506940 659104 511620 659704
rect 240858 657780 241818 658700
rect 329040 658684 329242 659104
rect 329040 658502 329240 658684
rect 329100 657980 329240 658502
rect 419260 658224 419460 659104
rect 509040 658684 509242 659104
rect 509040 658502 509240 658684
rect 329100 657962 329158 657980
rect 329142 657946 329158 657962
rect 329192 657962 329240 657980
rect 329192 657946 329204 657962
rect 329142 657944 329204 657946
rect 329146 657940 329204 657944
rect 237138 657180 241818 657780
rect 327920 657884 328720 657924
rect 327920 657724 327980 657884
rect 328140 657864 328720 657884
rect 329108 657896 329154 657908
rect 329108 657864 329114 657896
rect 328140 657744 329114 657864
rect 328140 657724 328720 657744
rect 327920 657684 328720 657724
rect 329108 657720 329114 657744
rect 329148 657720 329154 657896
rect 329108 657708 329154 657720
rect 329196 657896 329242 657908
rect 329196 657720 329202 657896
rect 329236 657864 329242 657896
rect 330160 657884 330360 657904
rect 330160 657864 330180 657884
rect 329236 657744 330180 657864
rect 329236 657720 329242 657744
rect 329196 657708 329242 657720
rect 330160 657724 330180 657744
rect 330340 657724 330360 657884
rect 330160 657704 330360 657724
rect 417920 657884 418660 657924
rect 417920 657724 417980 657884
rect 418140 657724 418660 657884
rect 417920 657684 418660 657724
rect 329146 657670 329204 657676
rect 329146 657664 329158 657670
rect 329100 657636 329158 657664
rect 329192 657664 329204 657670
rect 329192 657636 329240 657664
rect 59548 656640 59748 657180
rect 149238 656760 149440 657180
rect 59598 656061 59698 656640
rect 149238 656578 149438 656760
rect 59598 656055 59707 656061
rect 59598 656040 59627 656055
rect 59615 656021 59627 656040
rect 59695 656021 59707 656055
rect 149298 656056 149438 656578
rect 239258 656320 239498 657180
rect 329100 657124 329240 657636
rect 418460 657464 418660 657684
rect 419320 657547 419440 658224
rect 509100 657980 509240 658502
rect 509100 657962 509158 657980
rect 509142 657946 509158 657962
rect 509192 657962 509240 657980
rect 509192 657946 509204 657962
rect 509142 657944 509204 657946
rect 509146 657940 509204 657944
rect 419320 657513 419339 657547
rect 419407 657513 419440 657547
rect 419320 657504 419440 657513
rect 420160 657884 420360 657904
rect 420160 657724 420180 657884
rect 420340 657724 420360 657884
rect 419271 657464 419317 657466
rect 418460 657454 419317 657464
rect 418460 657278 419277 657454
rect 419311 657278 419317 657454
rect 418460 657266 419317 657278
rect 419429 657464 419475 657466
rect 420160 657464 420360 657724
rect 507920 657884 508720 657924
rect 507920 657724 507980 657884
rect 508140 657864 508720 657884
rect 509108 657896 509154 657908
rect 509108 657864 509114 657896
rect 508140 657744 509114 657864
rect 508140 657724 508720 657744
rect 507920 657684 508720 657724
rect 509108 657720 509114 657744
rect 509148 657720 509154 657896
rect 509108 657708 509154 657720
rect 509196 657896 509242 657908
rect 509196 657720 509202 657896
rect 509236 657864 509242 657896
rect 510160 657884 510360 657904
rect 510160 657864 510180 657884
rect 509236 657744 510180 657864
rect 509236 657720 509242 657744
rect 509196 657708 509242 657720
rect 510160 657724 510180 657744
rect 510340 657724 510360 657884
rect 510160 657704 510360 657724
rect 509146 657670 509204 657676
rect 509146 657664 509158 657670
rect 419429 657454 420360 657464
rect 419429 657278 419435 657454
rect 419469 657278 420360 657454
rect 419429 657266 420360 657278
rect 418460 657264 419300 657266
rect 419440 657264 420360 657266
rect 509100 657636 509158 657664
rect 509192 657664 509204 657670
rect 509192 657636 509240 657664
rect 419327 657224 419419 657225
rect 149298 656038 149356 656056
rect 59615 656015 59707 656021
rect 149340 656022 149356 656038
rect 149390 656038 149438 656056
rect 149390 656022 149402 656038
rect 239338 656033 239378 656320
rect 329040 656164 329240 657124
rect 419320 657219 419420 657224
rect 419320 657185 419339 657219
rect 419407 657185 419420 657219
rect 419320 656764 419420 657185
rect 509100 657124 509240 657636
rect 419260 656164 419460 656764
rect 509040 656164 509240 657124
rect 149340 656020 149402 656022
rect 149344 656016 149402 656020
rect 239327 656027 239385 656033
rect 58118 655960 58918 656000
rect 58118 655800 58178 655960
rect 58338 655940 58918 655960
rect 59559 655971 59605 655983
rect 59559 655940 59565 655971
rect 58338 655840 59565 655940
rect 58338 655800 58918 655840
rect 58118 655760 58918 655800
rect 59559 655795 59565 655840
rect 59599 655795 59605 655971
rect 59559 655783 59605 655795
rect 59717 655971 59763 655983
rect 59717 655795 59723 655971
rect 59757 655940 59763 655971
rect 60348 655960 60548 655990
rect 60348 655940 60378 655960
rect 59757 655840 60378 655940
rect 59757 655795 59763 655840
rect 59717 655783 59763 655795
rect 60348 655800 60378 655840
rect 60538 655800 60548 655960
rect 60348 655790 60548 655800
rect 148118 655960 148918 656000
rect 148118 655800 148178 655960
rect 148338 655940 148918 655960
rect 149306 655972 149352 655984
rect 149306 655940 149312 655972
rect 148338 655820 149312 655940
rect 148338 655800 148918 655820
rect 148118 655760 148918 655800
rect 149306 655796 149312 655820
rect 149346 655796 149352 655972
rect 149306 655784 149352 655796
rect 149394 655972 149440 655984
rect 238118 655980 238558 656000
rect 239327 655993 239339 656027
rect 239373 655993 239385 656027
rect 239327 655987 239385 655993
rect 149394 655796 149400 655972
rect 149434 655940 149440 655972
rect 150358 655960 150558 655980
rect 150358 655940 150378 655960
rect 149434 655820 150378 655940
rect 149434 655796 149440 655820
rect 149394 655784 149440 655796
rect 150358 655800 150378 655820
rect 150538 655800 150558 655960
rect 150358 655780 150558 655800
rect 238118 655960 238918 655980
rect 238118 655800 238178 655960
rect 238338 655900 238918 655960
rect 240078 655960 240558 655980
rect 239289 655934 239335 655946
rect 239289 655900 239295 655934
rect 238338 655840 239295 655900
rect 238338 655800 238918 655840
rect 238118 655760 238918 655800
rect 239289 655758 239295 655840
rect 239329 655758 239335 655934
rect 59615 655745 59707 655751
rect 59615 655740 59627 655745
rect 59598 655711 59627 655740
rect 59695 655711 59707 655745
rect 149344 655746 149402 655752
rect 239289 655746 239335 655758
rect 239377 655934 239423 655946
rect 239377 655758 239383 655934
rect 239417 655900 239423 655934
rect 240078 655900 240378 655960
rect 239417 655840 240378 655900
rect 239417 655758 239423 655840
rect 240078 655800 240378 655840
rect 240538 655800 240558 655960
rect 240078 655780 240558 655800
rect 239377 655746 239423 655758
rect 149344 655740 149356 655746
rect 59598 655705 59707 655711
rect 149298 655712 149356 655740
rect 149390 655740 149402 655746
rect 149390 655712 149438 655740
rect 59598 655290 59698 655705
rect 59548 654240 59748 655290
rect 149298 655200 149438 655712
rect 239327 655699 239385 655705
rect 239327 655665 239339 655699
rect 239373 655665 239385 655699
rect 239327 655659 239385 655665
rect 239338 655380 239378 655659
rect 326880 655564 331560 656164
rect 149238 654240 149438 655200
rect 239278 654240 239498 655380
rect 326880 654644 327840 655564
rect 57078 653640 61758 654240
rect 57078 652720 58038 653640
rect 57078 652120 57238 652720
rect 57838 652120 58038 652720
rect 57078 651960 58038 652120
rect 60798 652720 61758 653640
rect 60798 652120 60958 652720
rect 61558 652120 61758 652720
rect 60798 651960 61758 652120
rect 147078 653640 151758 654240
rect 147078 652720 148038 653640
rect 147078 652120 147238 652720
rect 147838 652120 148038 652720
rect 147078 651960 148038 652120
rect 150798 652720 151758 653640
rect 150798 652120 150958 652720
rect 151558 652120 151758 652720
rect 150798 651960 151758 652120
rect 237078 653640 241758 654240
rect 326880 654044 327040 654644
rect 327640 654044 327840 654644
rect 326880 653884 327840 654044
rect 330600 654644 331560 655564
rect 330600 654044 330760 654644
rect 331360 654044 331560 654644
rect 330600 653884 331560 654044
rect 416880 655564 421560 656164
rect 416880 654644 417840 655564
rect 416880 654044 417040 654644
rect 417640 654044 417840 654644
rect 416880 653884 417840 654044
rect 420600 654644 421560 655564
rect 420600 654044 420760 654644
rect 421360 654044 421560 654644
rect 420600 653884 421560 654044
rect 506880 655564 511560 656164
rect 506880 654644 507840 655564
rect 506880 654044 507040 654644
rect 507640 654044 507840 654644
rect 506880 653884 507840 654044
rect 510600 654644 511560 655564
rect 510600 654044 510760 654644
rect 511360 654044 511560 654644
rect 510600 653884 511560 654044
rect 237078 652720 238038 653640
rect 237078 652120 237238 652720
rect 237838 652120 238038 652720
rect 237078 651960 238038 652120
rect 240798 652720 241758 653640
rect 240798 652120 240958 652720
rect 241558 652120 241758 652720
rect 240798 651960 241758 652120
rect 416940 586224 417900 586384
rect 416940 585624 417100 586224
rect 417700 585624 417900 586224
rect 416940 584704 417900 585624
rect 420660 586224 421620 586384
rect 420660 585624 420820 586224
rect 421420 585624 421620 586224
rect 419000 584704 419300 584714
rect 420660 584704 421620 585624
rect 57138 584300 58098 584460
rect 57138 583700 57298 584300
rect 57898 583700 58098 584300
rect 57138 582780 58098 583700
rect 60858 584300 61818 584460
rect 60858 583700 61018 584300
rect 61618 583700 61818 584300
rect 59198 582780 59498 582790
rect 60858 582780 61818 583700
rect 57138 582190 61818 582780
rect 57138 582180 59238 582190
rect 59498 582180 61818 582190
rect 147138 584300 148098 584460
rect 147138 583700 147298 584300
rect 147898 583700 148098 584300
rect 147138 582780 148098 583700
rect 150858 584300 151818 584460
rect 150858 583700 151018 584300
rect 151618 583700 151818 584300
rect 150858 582780 151818 583700
rect 147138 582180 151818 582780
rect 237138 584300 238098 584460
rect 237138 583700 237298 584300
rect 237898 583700 238098 584300
rect 237138 582780 238098 583700
rect 240858 584300 241818 584460
rect 240858 583700 241018 584300
rect 241618 583700 241818 584300
rect 240858 582780 241818 583700
rect 237138 582180 241818 582780
rect 327138 584300 328098 584460
rect 327138 583700 327298 584300
rect 327898 583700 328098 584300
rect 327138 582780 328098 583700
rect 330858 584300 331818 584460
rect 330858 583700 331018 584300
rect 331618 583700 331818 584300
rect 416940 584114 421620 584704
rect 416940 584104 419040 584114
rect 419300 584104 421620 584114
rect 506940 586224 507900 586384
rect 506940 585624 507100 586224
rect 507700 585624 507900 586224
rect 506940 584704 507900 585624
rect 510660 586224 511620 586384
rect 510660 585624 510820 586224
rect 511420 585624 511620 586224
rect 510660 584704 511620 585624
rect 506940 584104 511620 584704
rect 330858 582780 331818 583700
rect 419350 583564 419550 584104
rect 419400 582985 419500 583564
rect 509360 583444 509580 584104
rect 419400 582979 419509 582985
rect 419400 582964 419429 582979
rect 419417 582945 419429 582964
rect 419497 582945 419509 582979
rect 419417 582939 419509 582945
rect 327138 582180 331818 582780
rect 417920 582884 418720 582924
rect 417920 582724 417980 582884
rect 418140 582864 418720 582884
rect 419361 582895 419407 582907
rect 419361 582864 419367 582895
rect 418140 582764 419367 582864
rect 418140 582724 418720 582764
rect 417920 582684 418720 582724
rect 419361 582719 419367 582764
rect 419401 582719 419407 582895
rect 419361 582707 419407 582719
rect 419519 582895 419565 582907
rect 419519 582719 419525 582895
rect 419559 582864 419565 582895
rect 420150 582884 420350 582914
rect 420150 582864 420180 582884
rect 419559 582764 420180 582864
rect 419559 582719 419565 582764
rect 419519 582707 419565 582719
rect 420150 582724 420180 582764
rect 420340 582724 420350 582884
rect 420150 582714 420350 582724
rect 507920 582884 508660 582924
rect 507920 582724 507980 582884
rect 508140 582724 508660 582884
rect 507920 582684 508660 582724
rect 419417 582669 419509 582675
rect 419417 582664 419429 582669
rect 419400 582635 419429 582664
rect 419497 582635 419509 582669
rect 419400 582629 419509 582635
rect 419400 582214 419500 582629
rect 508460 582584 508660 582684
rect 509420 582689 509520 583444
rect 509420 582664 509439 582689
rect 509427 582655 509439 582664
rect 509507 582664 509520 582689
rect 510160 582884 510360 582904
rect 510160 582724 510180 582884
rect 510340 582724 510360 582884
rect 509507 582655 509519 582664
rect 509427 582649 509519 582655
rect 509371 582605 509417 582617
rect 509371 582584 509377 582605
rect 508460 582484 509377 582584
rect 508460 582424 508660 582484
rect 509371 582429 509377 582484
rect 509411 582429 509417 582605
rect 509371 582417 509417 582429
rect 509529 582605 509575 582617
rect 509529 582429 509535 582605
rect 509569 582584 509575 582605
rect 510160 582584 510360 582724
rect 509569 582484 510360 582584
rect 509569 582429 509575 582484
rect 509529 582417 509575 582429
rect 510160 582424 510360 582484
rect 509427 582384 509519 582385
rect 509420 582379 509519 582384
rect 509420 582345 509439 582379
rect 509507 582345 509519 582379
rect 509420 582339 509519 582345
rect 59548 581640 59748 582180
rect 59598 581061 59698 581640
rect 149558 581520 149778 582180
rect 239238 581760 239440 582180
rect 239238 581578 239438 581760
rect 59598 581055 59707 581061
rect 59598 581040 59627 581055
rect 59615 581021 59627 581040
rect 59695 581021 59707 581055
rect 59615 581015 59707 581021
rect 58118 580960 58918 581000
rect 58118 580800 58178 580960
rect 58338 580940 58918 580960
rect 59559 580971 59605 580983
rect 59559 580940 59565 580971
rect 58338 580840 59565 580940
rect 58338 580800 58918 580840
rect 58118 580760 58918 580800
rect 59559 580795 59565 580840
rect 59599 580795 59605 580971
rect 59559 580783 59605 580795
rect 59717 580971 59763 580983
rect 59717 580795 59723 580971
rect 59757 580940 59763 580971
rect 60348 580960 60548 580990
rect 60348 580940 60378 580960
rect 59757 580840 60378 580940
rect 59757 580795 59763 580840
rect 59717 580783 59763 580795
rect 60348 580800 60378 580840
rect 60538 580800 60548 580960
rect 60348 580790 60548 580800
rect 148118 580960 148858 581000
rect 148118 580800 148178 580960
rect 148338 580800 148858 580960
rect 148118 580760 148858 580800
rect 59615 580745 59707 580751
rect 59615 580740 59627 580745
rect 59598 580711 59627 580740
rect 59695 580711 59707 580745
rect 59598 580705 59707 580711
rect 59598 580290 59698 580705
rect 148658 580660 148858 580760
rect 149618 580765 149718 581520
rect 239298 581056 239438 581578
rect 329458 581300 329658 582180
rect 239298 581038 239356 581056
rect 239340 581022 239356 581038
rect 239390 581038 239438 581056
rect 239390 581022 239402 581038
rect 239340 581020 239402 581022
rect 239344 581016 239402 581020
rect 149618 580740 149637 580765
rect 149625 580731 149637 580740
rect 149705 580740 149718 580765
rect 150358 580960 150558 580980
rect 150358 580800 150378 580960
rect 150538 580800 150558 580960
rect 149705 580731 149717 580740
rect 149625 580725 149717 580731
rect 149569 580681 149615 580693
rect 149569 580660 149575 580681
rect 148658 580560 149575 580660
rect 148658 580500 148858 580560
rect 149569 580505 149575 580560
rect 149609 580505 149615 580681
rect 149569 580493 149615 580505
rect 149727 580681 149773 580693
rect 149727 580505 149733 580681
rect 149767 580660 149773 580681
rect 150358 580660 150558 580800
rect 238118 580960 238918 581000
rect 238118 580800 238178 580960
rect 238338 580940 238918 580960
rect 239306 580972 239352 580984
rect 239306 580940 239312 580972
rect 238338 580820 239312 580940
rect 238338 580800 238918 580820
rect 238118 580760 238918 580800
rect 239306 580796 239312 580820
rect 239346 580796 239352 580972
rect 239306 580784 239352 580796
rect 239394 580972 239440 580984
rect 239394 580796 239400 580972
rect 239434 580940 239440 580972
rect 240358 580960 240558 580980
rect 240358 580940 240378 580960
rect 239434 580820 240378 580940
rect 239434 580796 239440 580820
rect 239394 580784 239440 580796
rect 240358 580800 240378 580820
rect 240538 580800 240558 580960
rect 240358 580780 240558 580800
rect 328118 580960 328858 581000
rect 328118 580800 328178 580960
rect 328338 580800 328858 580960
rect 328118 580760 328858 580800
rect 239344 580746 239402 580752
rect 239344 580740 239356 580746
rect 149767 580560 150558 580660
rect 149767 580505 149773 580560
rect 149727 580493 149773 580505
rect 150358 580500 150558 580560
rect 239298 580712 239356 580740
rect 239390 580740 239402 580746
rect 239390 580712 239438 580740
rect 149625 580460 149717 580461
rect 149618 580455 149717 580460
rect 149618 580421 149637 580455
rect 149705 580421 149717 580455
rect 149618 580415 149717 580421
rect 59548 579240 59748 580290
rect 149618 579900 149698 580415
rect 239298 580200 239438 580712
rect 328658 580540 328858 580760
rect 329518 580623 329638 581300
rect 419350 581164 419550 582214
rect 509420 581824 509500 582339
rect 509360 581164 509560 581824
rect 329518 580589 329537 580623
rect 329605 580589 329638 580623
rect 329518 580580 329638 580589
rect 330358 580960 330558 580980
rect 330358 580800 330378 580960
rect 330538 580800 330558 580960
rect 329469 580540 329515 580542
rect 328658 580530 329515 580540
rect 328658 580354 329475 580530
rect 329509 580354 329515 580530
rect 328658 580342 329515 580354
rect 329627 580540 329673 580542
rect 330358 580540 330558 580800
rect 329627 580530 330558 580540
rect 329627 580354 329633 580530
rect 329667 580354 330558 580530
rect 329627 580342 330558 580354
rect 328658 580340 329498 580342
rect 329638 580340 330558 580342
rect 416880 580564 421560 581164
rect 329525 580300 329617 580301
rect 149558 579240 149758 579900
rect 239238 579240 239438 580200
rect 329518 580295 329618 580300
rect 329518 580261 329537 580295
rect 329605 580261 329618 580295
rect 329518 579840 329618 580261
rect 329458 579240 329658 579840
rect 416880 579644 417840 580564
rect 57078 578640 61758 579240
rect 57078 577720 58038 578640
rect 57078 577120 57238 577720
rect 57838 577120 58038 577720
rect 57078 576960 58038 577120
rect 60798 577720 61758 578640
rect 60798 577120 60958 577720
rect 61558 577120 61758 577720
rect 60798 576960 61758 577120
rect 147078 578640 151758 579240
rect 147078 577720 148038 578640
rect 147078 577120 147238 577720
rect 147838 577120 148038 577720
rect 147078 576960 148038 577120
rect 150798 577720 151758 578640
rect 150798 577120 150958 577720
rect 151558 577120 151758 577720
rect 150798 576960 151758 577120
rect 237078 578640 241758 579240
rect 237078 577720 238038 578640
rect 237078 577120 237238 577720
rect 237838 577120 238038 577720
rect 237078 576960 238038 577120
rect 240798 577720 241758 578640
rect 240798 577120 240958 577720
rect 241558 577120 241758 577720
rect 240798 576960 241758 577120
rect 327078 578640 331758 579240
rect 416880 579044 417040 579644
rect 417640 579044 417840 579644
rect 416880 578884 417840 579044
rect 420600 579644 421560 580564
rect 420600 579044 420760 579644
rect 421360 579044 421560 579644
rect 420600 578884 421560 579044
rect 506880 580564 511560 581164
rect 506880 579644 507840 580564
rect 506880 579044 507040 579644
rect 507640 579044 507840 579644
rect 506880 578884 507840 579044
rect 510600 579644 511560 580564
rect 510600 579044 510760 579644
rect 511360 579044 511560 579644
rect 510600 578884 511560 579044
rect 327078 577720 328038 578640
rect 327078 577120 327238 577720
rect 327838 577120 328038 577720
rect 327078 576960 328038 577120
rect 330798 577720 331758 578640
rect 330798 577120 330958 577720
rect 331558 577120 331758 577720
rect 330798 576960 331758 577120
rect 64394 504794 65846 505158
rect 64394 503970 64790 504794
rect 65516 503970 65846 504794
rect 57138 495400 58098 495560
rect 57138 494800 57298 495400
rect 57898 494800 58098 495400
rect 57138 493880 58098 494800
rect 60858 495400 61818 495560
rect 60858 494800 61018 495400
rect 61618 494800 61818 495400
rect 64394 494824 65846 503970
rect 154394 504794 155846 505158
rect 154394 503970 154790 504794
rect 155516 503970 155846 504794
rect 154394 498735 155846 503970
rect 244394 504794 245846 505158
rect 244394 503970 244790 504794
rect 245516 503970 245846 504794
rect 244394 495113 245846 503970
rect 334394 504794 335846 505158
rect 334394 503970 334790 504794
rect 335516 503970 335846 504794
rect 334394 494824 335846 503970
rect 424394 504794 425846 505158
rect 424394 503970 424790 504794
rect 425516 503970 425846 504794
rect 417138 495400 418098 495560
rect 60858 493880 61818 494800
rect 57138 493280 61818 493880
rect 417138 494800 417298 495400
rect 417898 494800 418098 495400
rect 417138 493880 418098 494800
rect 420858 495400 421818 495560
rect 420858 494800 421018 495400
rect 421618 494800 421818 495400
rect 424394 494824 425846 503970
rect 514394 504794 515846 505158
rect 514394 503970 514790 504794
rect 515516 503970 515846 504794
rect 507138 495400 508098 495560
rect 420858 493880 421818 494800
rect 323744 493502 324264 493736
rect 323744 493378 323908 493502
rect 324016 493378 324264 493502
rect 59380 492678 59564 493280
rect 230433 492790 231381 492796
rect 59368 492592 60088 492678
rect 60002 492392 60088 492592
rect 60002 492328 60008 492392
rect 60080 492328 60088 492392
rect 60002 492302 60088 492328
rect 59006 491996 62804 492050
rect 58891 491843 58983 491849
rect 57964 491786 58164 491834
rect 58891 491809 58903 491843
rect 58971 491809 58983 491843
rect 58891 491803 58983 491809
rect 57964 491684 57996 491786
rect 58146 491684 58164 491786
rect 57964 491634 58164 491684
rect 58828 491771 58860 491788
rect 59012 491771 59042 491996
rect 58828 491759 58881 491771
rect 58828 491699 58841 491759
rect 58875 491699 58881 491759
rect 58828 491687 58881 491699
rect 58993 491759 59042 491771
rect 58993 491699 58999 491759
rect 59033 491699 59042 491759
rect 58993 491687 59042 491699
rect 58039 491434 58085 491634
rect 58828 491434 58860 491687
rect 59012 491666 59042 491687
rect 59102 491771 59132 491996
rect 59167 491843 59259 491849
rect 59167 491809 59179 491843
rect 59247 491809 59259 491843
rect 59167 491803 59259 491809
rect 59443 491843 59535 491849
rect 59443 491809 59455 491843
rect 59523 491809 59535 491843
rect 59443 491803 59535 491809
rect 59294 491771 59326 491790
rect 59102 491759 59157 491771
rect 59102 491699 59117 491759
rect 59151 491699 59157 491759
rect 59102 491687 59157 491699
rect 59269 491759 59326 491771
rect 59269 491699 59275 491759
rect 59309 491699 59326 491759
rect 59269 491687 59326 491699
rect 59102 491666 59132 491687
rect 58891 491649 58983 491655
rect 58891 491615 58903 491649
rect 58971 491615 58983 491649
rect 58891 491609 58983 491615
rect 59167 491649 59259 491655
rect 59167 491615 59179 491649
rect 59247 491615 59259 491649
rect 59167 491609 59259 491615
rect 59294 491434 59326 491687
rect 59376 491771 59408 491790
rect 59564 491771 59594 491996
rect 59376 491759 59433 491771
rect 59376 491699 59393 491759
rect 59427 491699 59433 491759
rect 59376 491687 59433 491699
rect 59545 491759 59594 491771
rect 59545 491699 59551 491759
rect 59585 491699 59594 491759
rect 59545 491687 59594 491699
rect 59376 491434 59408 491687
rect 59564 491668 59594 491687
rect 59654 491771 59684 491996
rect 60006 491872 60086 491882
rect 60006 491849 60008 491872
rect 59719 491843 59811 491849
rect 59719 491809 59731 491843
rect 59799 491809 59811 491843
rect 59719 491803 59811 491809
rect 59995 491843 60008 491849
rect 60076 491849 60086 491872
rect 59995 491809 60007 491843
rect 60076 491816 60087 491849
rect 60075 491809 60087 491816
rect 59995 491803 60087 491809
rect 59846 491771 59878 491790
rect 59654 491759 59709 491771
rect 59654 491699 59669 491759
rect 59703 491699 59709 491759
rect 59654 491687 59709 491699
rect 59821 491759 59878 491771
rect 59821 491699 59827 491759
rect 59861 491699 59878 491759
rect 59821 491687 59878 491699
rect 59654 491666 59684 491687
rect 59443 491649 59535 491655
rect 59443 491615 59455 491649
rect 59523 491615 59535 491649
rect 59443 491609 59535 491615
rect 59719 491649 59811 491655
rect 59719 491615 59731 491649
rect 59799 491615 59811 491649
rect 59719 491609 59811 491615
rect 59846 491434 59878 491687
rect 59934 491771 59966 491788
rect 60118 491771 60148 491996
rect 59934 491759 59985 491771
rect 59934 491699 59945 491759
rect 59979 491699 59985 491759
rect 59934 491687 59985 491699
rect 60097 491759 60148 491771
rect 60097 491699 60103 491759
rect 60137 491699 60148 491759
rect 60097 491687 60148 491699
rect 59934 491434 59966 491687
rect 60118 491662 60148 491687
rect 60208 491771 60238 491996
rect 60271 491843 60363 491849
rect 60271 491809 60283 491843
rect 60351 491809 60363 491843
rect 60271 491803 60363 491809
rect 60547 491843 60639 491849
rect 60547 491809 60559 491843
rect 60627 491809 60639 491843
rect 60547 491803 60639 491809
rect 60394 491771 60426 491790
rect 60208 491759 60261 491771
rect 60208 491699 60221 491759
rect 60255 491699 60261 491759
rect 60208 491687 60261 491699
rect 60373 491759 60426 491771
rect 60373 491699 60379 491759
rect 60413 491699 60426 491759
rect 60373 491687 60426 491699
rect 60208 491660 60238 491687
rect 60000 491655 60080 491656
rect 59995 491649 60087 491655
rect 59995 491615 60007 491649
rect 60075 491642 60087 491649
rect 59995 491609 60008 491615
rect 60000 491586 60008 491609
rect 60076 491609 60087 491642
rect 60271 491649 60363 491655
rect 60271 491615 60283 491649
rect 60351 491615 60363 491649
rect 60271 491609 60363 491615
rect 60076 491586 60080 491609
rect 60000 491578 60080 491586
rect 60394 491434 60426 491687
rect 60482 491771 60514 491788
rect 60668 491771 60698 491996
rect 60482 491759 60537 491771
rect 60482 491699 60497 491759
rect 60531 491699 60537 491759
rect 60482 491687 60537 491699
rect 60649 491759 60698 491771
rect 60649 491699 60655 491759
rect 60689 491699 60698 491759
rect 60649 491687 60698 491699
rect 60482 491434 60514 491687
rect 60668 491672 60698 491687
rect 60758 491771 60788 491996
rect 60823 491843 60915 491849
rect 60823 491809 60835 491843
rect 60903 491809 60915 491843
rect 60823 491803 60915 491809
rect 61099 491843 61191 491849
rect 61099 491809 61111 491843
rect 61179 491809 61191 491843
rect 61099 491803 61191 491809
rect 60946 491771 60978 491790
rect 60758 491759 60813 491771
rect 60758 491699 60773 491759
rect 60807 491699 60813 491759
rect 60758 491687 60813 491699
rect 60925 491759 60978 491771
rect 60925 491699 60931 491759
rect 60965 491699 60978 491759
rect 60925 491687 60978 491699
rect 60758 491672 60788 491687
rect 60547 491649 60639 491655
rect 60547 491615 60559 491649
rect 60627 491615 60639 491649
rect 60547 491609 60639 491615
rect 60823 491649 60915 491655
rect 60823 491615 60835 491649
rect 60903 491615 60915 491649
rect 60823 491609 60915 491615
rect 60946 491434 60978 491687
rect 61030 491771 61062 491782
rect 61222 491771 61252 491996
rect 61030 491759 61089 491771
rect 61030 491699 61049 491759
rect 61083 491699 61089 491759
rect 61030 491687 61089 491699
rect 61201 491759 61252 491771
rect 61201 491699 61207 491759
rect 61241 491699 61252 491759
rect 61201 491687 61252 491699
rect 61030 491434 61062 491687
rect 61222 491672 61252 491687
rect 61306 491771 61336 491996
rect 61375 491843 61467 491849
rect 61375 491809 61387 491843
rect 61455 491809 61467 491843
rect 61375 491803 61467 491809
rect 61496 491771 61528 491790
rect 61306 491759 61365 491771
rect 61306 491699 61325 491759
rect 61359 491699 61365 491759
rect 61306 491687 61365 491699
rect 61477 491759 61528 491771
rect 61477 491699 61483 491759
rect 61517 491699 61528 491759
rect 61477 491687 61528 491699
rect 61306 491674 61336 491687
rect 61099 491649 61191 491655
rect 61099 491615 61111 491649
rect 61179 491615 61191 491649
rect 61099 491609 61191 491615
rect 61375 491649 61467 491655
rect 61375 491615 61387 491649
rect 61455 491615 61467 491649
rect 61375 491609 61467 491615
rect 61496 491434 61528 491687
rect 61620 491576 61658 491996
rect 62747 491818 62801 491996
rect 62668 491786 62868 491818
rect 62668 491638 62696 491786
rect 62844 491638 62868 491786
rect 62668 491618 62868 491638
rect 141258 491469 142348 492005
rect 323744 492700 324264 493378
rect 417138 493280 421818 493880
rect 507138 494800 507298 495400
rect 507898 494800 508098 495400
rect 507138 493880 508098 494800
rect 510858 495400 511818 495560
rect 510858 494800 511018 495400
rect 511618 494800 511818 495400
rect 514394 494824 515846 503970
rect 510858 493880 511818 494800
rect 507138 493280 511818 493880
rect 323888 492598 323972 492700
rect 323888 492556 323904 492598
rect 323958 492556 323972 492598
rect 323888 492536 323972 492556
rect 338790 492400 339590 492534
rect 321787 492028 321793 492354
rect 322119 492146 322656 492354
rect 324001 492334 339590 492400
rect 323881 492231 323973 492237
rect 323881 492197 323893 492231
rect 323961 492197 323973 492231
rect 323881 492191 323973 492197
rect 324006 492159 324046 492334
rect 323825 492147 323871 492159
rect 323825 492146 323831 492147
rect 322119 492088 323831 492146
rect 322119 492028 322656 492088
rect 323667 491910 323709 492088
rect 323825 492087 323831 492088
rect 323865 492087 323871 492147
rect 323825 492075 323871 492087
rect 323983 492147 324046 492159
rect 323983 492087 323989 492147
rect 324023 492087 324046 492147
rect 323983 492075 324046 492087
rect 324006 492068 324046 492075
rect 324088 492159 324128 492334
rect 324157 492231 324249 492237
rect 324157 492197 324169 492231
rect 324237 492197 324249 492231
rect 324157 492191 324249 492197
rect 324433 492231 324525 492237
rect 324433 492197 324445 492231
rect 324513 492197 324525 492231
rect 324433 492191 324525 492197
rect 324282 492159 324312 492166
rect 324088 492147 324147 492159
rect 324088 492087 324107 492147
rect 324141 492087 324147 492147
rect 324088 492075 324147 492087
rect 324259 492147 324312 492159
rect 324259 492087 324265 492147
rect 324299 492087 324312 492147
rect 324259 492075 324312 492087
rect 324088 492070 324128 492075
rect 323881 492037 323973 492043
rect 323881 492003 323893 492037
rect 323961 492003 323973 492037
rect 323881 491997 323973 492003
rect 324157 492037 324249 492043
rect 324157 492003 324169 492037
rect 324237 492003 324249 492037
rect 324157 491997 324249 492003
rect 323839 491910 324015 491911
rect 324282 491910 324312 492075
rect 324368 492159 324398 492166
rect 324564 492159 324604 492334
rect 324368 492147 324423 492159
rect 324368 492087 324383 492147
rect 324417 492087 324423 492147
rect 324368 492075 324423 492087
rect 324535 492147 324604 492159
rect 324535 492087 324541 492147
rect 324575 492087 324604 492147
rect 324535 492075 324604 492087
rect 324368 491910 324398 492075
rect 324564 492070 324604 492075
rect 324632 492159 324672 492334
rect 324709 492231 324801 492237
rect 324709 492197 324721 492231
rect 324789 492197 324801 492231
rect 324709 492191 324801 492197
rect 324985 492231 325077 492237
rect 324985 492197 324997 492231
rect 325065 492197 325077 492231
rect 324985 492191 325077 492197
rect 324836 492159 324866 492166
rect 324632 492147 324699 492159
rect 324632 492087 324659 492147
rect 324693 492087 324699 492147
rect 324632 492075 324699 492087
rect 324811 492147 324866 492159
rect 324811 492087 324817 492147
rect 324851 492087 324866 492147
rect 324811 492075 324866 492087
rect 324632 492070 324672 492075
rect 324433 492037 324525 492043
rect 324433 492003 324445 492037
rect 324513 492003 324525 492037
rect 324433 491997 324525 492003
rect 324709 492037 324801 492043
rect 324709 492003 324721 492037
rect 324789 492003 324801 492037
rect 324709 491997 324801 492003
rect 324836 491910 324866 492075
rect 324922 492159 324952 492166
rect 325112 492159 325152 492334
rect 324922 492147 324975 492159
rect 324922 492087 324935 492147
rect 324969 492087 324975 492147
rect 324922 492075 324975 492087
rect 325087 492147 325152 492159
rect 325087 492087 325093 492147
rect 325127 492087 325152 492147
rect 325087 492075 325152 492087
rect 324922 491910 324952 492075
rect 325112 492066 325152 492075
rect 325184 492159 325224 492334
rect 325261 492231 325353 492237
rect 325261 492197 325273 492231
rect 325341 492197 325353 492231
rect 325261 492191 325353 492197
rect 325537 492231 325629 492237
rect 325537 492197 325549 492231
rect 325617 492197 325629 492231
rect 325537 492191 325629 492197
rect 325384 492159 325414 492166
rect 325184 492147 325251 492159
rect 325184 492087 325211 492147
rect 325245 492087 325251 492147
rect 325184 492075 325251 492087
rect 325363 492147 325414 492159
rect 325363 492087 325369 492147
rect 325403 492087 325414 492147
rect 325363 492075 325414 492087
rect 325184 492070 325224 492075
rect 324985 492037 325077 492043
rect 324985 492003 324997 492037
rect 325065 492003 325077 492037
rect 324985 491997 325077 492003
rect 325261 492037 325353 492043
rect 325261 492003 325273 492037
rect 325341 492003 325353 492037
rect 325261 491997 325353 492003
rect 325384 491910 325414 492075
rect 325476 492159 325506 492164
rect 325664 492159 325704 492334
rect 325476 492147 325527 492159
rect 325476 492087 325487 492147
rect 325521 492087 325527 492147
rect 325476 492075 325527 492087
rect 325639 492147 325704 492159
rect 325639 492087 325645 492147
rect 325679 492087 325704 492147
rect 325639 492075 325704 492087
rect 325476 491910 325506 492075
rect 325664 492074 325704 492075
rect 325744 492159 325784 492334
rect 325813 492231 325905 492237
rect 325813 492197 325825 492231
rect 325893 492197 325905 492231
rect 325813 492191 325905 492197
rect 326089 492231 326181 492237
rect 326089 492197 326101 492231
rect 326169 492197 326181 492231
rect 326089 492191 326181 492197
rect 325934 492159 325964 492164
rect 325744 492147 325803 492159
rect 325744 492087 325763 492147
rect 325797 492087 325803 492147
rect 325744 492075 325803 492087
rect 325915 492147 325964 492159
rect 325915 492087 325921 492147
rect 325955 492087 325964 492147
rect 325915 492075 325964 492087
rect 325744 492074 325784 492075
rect 325537 492037 325629 492043
rect 325537 492003 325549 492037
rect 325617 492003 325629 492037
rect 325537 491997 325629 492003
rect 325813 492037 325905 492043
rect 325813 492003 325825 492037
rect 325893 492003 325905 492037
rect 325813 491997 325905 492003
rect 325934 491910 325964 492075
rect 326026 492159 326056 492162
rect 326218 492159 326258 492334
rect 326026 492147 326079 492159
rect 326026 492087 326039 492147
rect 326073 492087 326079 492147
rect 326026 492075 326079 492087
rect 326191 492147 326258 492159
rect 326191 492087 326197 492147
rect 326231 492087 326258 492147
rect 326191 492075 326258 492087
rect 326026 491910 326056 492075
rect 326218 492070 326258 492075
rect 326292 492159 326332 492334
rect 326365 492231 326457 492237
rect 326365 492197 326377 492231
rect 326445 492197 326457 492231
rect 326365 492191 326457 492197
rect 326641 492231 326733 492237
rect 326641 492197 326653 492231
rect 326721 492197 326733 492231
rect 326641 492191 326733 492197
rect 326490 492159 326520 492162
rect 326292 492147 326355 492159
rect 326292 492087 326315 492147
rect 326349 492087 326355 492147
rect 326292 492075 326355 492087
rect 326467 492147 326520 492159
rect 326467 492087 326473 492147
rect 326507 492087 326520 492147
rect 326467 492075 326520 492087
rect 326292 492072 326332 492075
rect 326089 492037 326181 492043
rect 326089 492003 326101 492037
rect 326169 492003 326181 492037
rect 326089 491997 326181 492003
rect 326365 492037 326457 492043
rect 326365 492003 326377 492037
rect 326445 492003 326457 492037
rect 326365 491997 326457 492003
rect 326490 491910 326520 492075
rect 326578 492159 326608 492160
rect 326770 492159 326810 492334
rect 326578 492147 326631 492159
rect 326578 492087 326591 492147
rect 326625 492087 326631 492147
rect 326578 492075 326631 492087
rect 326743 492147 326810 492159
rect 326743 492087 326749 492147
rect 326783 492087 326810 492147
rect 326743 492075 326810 492087
rect 326578 491910 326608 492075
rect 326770 492068 326810 492075
rect 326840 492159 326880 492334
rect 326917 492231 327009 492237
rect 326917 492197 326929 492231
rect 326997 492197 327009 492231
rect 326917 492191 327009 492197
rect 327193 492231 327285 492237
rect 327193 492197 327205 492231
rect 327273 492197 327285 492231
rect 327193 492191 327285 492197
rect 327040 492159 327070 492160
rect 326840 492147 326907 492159
rect 326840 492087 326867 492147
rect 326901 492087 326907 492147
rect 326840 492075 326907 492087
rect 327019 492147 327070 492159
rect 327019 492087 327025 492147
rect 327059 492087 327070 492147
rect 327019 492075 327070 492087
rect 326840 492072 326880 492075
rect 326641 492037 326733 492043
rect 326641 492003 326653 492037
rect 326721 492003 326733 492037
rect 326641 491997 326733 492003
rect 326917 492037 327009 492043
rect 326917 492003 326929 492037
rect 326997 492003 327009 492037
rect 326917 491997 327009 492003
rect 327040 491910 327070 492075
rect 327128 492159 327158 492160
rect 327318 492159 327358 492334
rect 327128 492147 327183 492159
rect 327128 492087 327143 492147
rect 327177 492087 327183 492147
rect 327128 492075 327183 492087
rect 327295 492147 327358 492159
rect 327295 492087 327301 492147
rect 327335 492087 327358 492147
rect 327295 492075 327358 492087
rect 327128 491910 327158 492075
rect 327318 492068 327358 492075
rect 327396 492159 327436 492334
rect 327469 492231 327561 492237
rect 327469 492197 327481 492231
rect 327549 492197 327561 492231
rect 327469 492191 327561 492197
rect 327745 492231 327837 492237
rect 327745 492197 327757 492231
rect 327825 492197 327837 492231
rect 327745 492191 327837 492197
rect 327592 492159 327622 492162
rect 327396 492147 327459 492159
rect 327396 492087 327419 492147
rect 327453 492087 327459 492147
rect 327396 492075 327459 492087
rect 327571 492147 327622 492159
rect 327571 492087 327577 492147
rect 327611 492087 327622 492147
rect 327571 492075 327622 492087
rect 327396 492072 327436 492075
rect 327193 492037 327285 492043
rect 327193 492003 327205 492037
rect 327273 492003 327285 492037
rect 327193 491997 327285 492003
rect 327469 492037 327561 492043
rect 327469 492003 327481 492037
rect 327549 492003 327561 492037
rect 327469 491997 327561 492003
rect 327592 491910 327622 492075
rect 327680 492159 327710 492162
rect 327872 492159 327912 492334
rect 327680 492147 327735 492159
rect 327680 492087 327695 492147
rect 327729 492087 327735 492147
rect 327680 492075 327735 492087
rect 327847 492147 327912 492159
rect 327847 492087 327853 492147
rect 327887 492087 327912 492147
rect 327847 492075 327912 492087
rect 327680 491910 327710 492075
rect 327872 492060 327912 492075
rect 327950 492159 327990 492334
rect 328021 492231 328113 492237
rect 328021 492197 328033 492231
rect 328101 492197 328113 492231
rect 328021 492191 328113 492197
rect 328297 492231 328389 492237
rect 328297 492197 328309 492231
rect 328377 492197 328389 492231
rect 328297 492191 328389 492197
rect 328144 492159 328174 492162
rect 327950 492147 328011 492159
rect 327950 492087 327971 492147
rect 328005 492087 328011 492147
rect 327950 492075 328011 492087
rect 328123 492147 328174 492159
rect 328123 492087 328129 492147
rect 328163 492087 328174 492147
rect 328123 492075 328174 492087
rect 327950 492068 327990 492075
rect 327745 492037 327837 492043
rect 327745 492003 327757 492037
rect 327825 492003 327837 492037
rect 327745 491997 327837 492003
rect 328021 492037 328113 492043
rect 328021 492003 328033 492037
rect 328101 492003 328113 492037
rect 328021 491997 328113 492003
rect 328144 491910 328174 492075
rect 328236 492159 328266 492162
rect 328428 492159 328468 492334
rect 328236 492147 328287 492159
rect 328236 492087 328247 492147
rect 328281 492087 328287 492147
rect 328236 492075 328287 492087
rect 328399 492147 328468 492159
rect 328399 492087 328405 492147
rect 328439 492087 328468 492147
rect 328399 492075 328468 492087
rect 328236 491910 328266 492075
rect 328428 492070 328468 492075
rect 328502 492159 328542 492334
rect 328573 492231 328665 492237
rect 328573 492197 328585 492231
rect 328653 492197 328665 492231
rect 328573 492191 328665 492197
rect 328849 492231 328941 492237
rect 328849 492197 328861 492231
rect 328929 492197 328941 492231
rect 328849 492191 328941 492197
rect 328698 492159 328728 492172
rect 328502 492147 328563 492159
rect 328502 492087 328523 492147
rect 328557 492087 328563 492147
rect 328502 492075 328563 492087
rect 328675 492147 328728 492159
rect 328675 492087 328681 492147
rect 328715 492087 328728 492147
rect 328675 492075 328728 492087
rect 328502 492074 328542 492075
rect 328297 492037 328389 492043
rect 328297 492003 328309 492037
rect 328377 492003 328389 492037
rect 328297 491997 328389 492003
rect 328573 492037 328665 492043
rect 328573 492003 328585 492037
rect 328653 492003 328665 492037
rect 328573 491997 328665 492003
rect 328698 491910 328728 492075
rect 328784 492159 328814 492170
rect 328972 492159 329006 492334
rect 328784 492147 328839 492159
rect 328784 492087 328799 492147
rect 328833 492087 328839 492147
rect 328784 492075 328839 492087
rect 328951 492147 329006 492159
rect 328951 492087 328957 492147
rect 328991 492087 329006 492147
rect 328951 492075 329006 492087
rect 328784 491910 328814 492075
rect 328972 492070 329006 492075
rect 329062 492159 329096 492334
rect 329125 492231 329217 492237
rect 329125 492197 329137 492231
rect 329205 492197 329217 492231
rect 329125 492191 329217 492197
rect 329401 492231 329493 492237
rect 329401 492197 329413 492231
rect 329481 492197 329493 492231
rect 329401 492191 329493 492197
rect 329252 492159 329282 492168
rect 329062 492147 329115 492159
rect 329062 492087 329075 492147
rect 329109 492087 329115 492147
rect 329062 492075 329115 492087
rect 329227 492147 329282 492159
rect 329227 492087 329233 492147
rect 329267 492087 329282 492147
rect 329227 492075 329282 492087
rect 329062 492070 329096 492075
rect 328849 492037 328941 492043
rect 328849 492003 328861 492037
rect 328929 492003 328941 492037
rect 328849 491997 328941 492003
rect 329125 492037 329217 492043
rect 329125 492003 329137 492037
rect 329205 492003 329217 492037
rect 329125 491997 329217 492003
rect 329252 491910 329282 492075
rect 329338 492159 329368 492168
rect 329528 492159 329562 492334
rect 329338 492147 329391 492159
rect 329338 492087 329351 492147
rect 329385 492087 329391 492147
rect 329338 492075 329391 492087
rect 329503 492147 329562 492159
rect 329503 492087 329509 492147
rect 329543 492087 329562 492147
rect 329503 492075 329562 492087
rect 329338 491910 329368 492075
rect 329528 492070 329562 492075
rect 329612 492159 329646 492334
rect 329677 492231 329769 492237
rect 329677 492197 329689 492231
rect 329757 492197 329769 492231
rect 329677 492191 329769 492197
rect 329804 492159 329838 492172
rect 329612 492147 329667 492159
rect 329612 492087 329627 492147
rect 329661 492087 329667 492147
rect 329612 492075 329667 492087
rect 329779 492147 329838 492159
rect 329779 492087 329785 492147
rect 329819 492087 329838 492147
rect 329779 492075 329838 492087
rect 329612 492074 329646 492075
rect 329401 492037 329493 492043
rect 329401 492003 329413 492037
rect 329481 492003 329493 492037
rect 329401 491997 329493 492003
rect 329677 492037 329769 492043
rect 329677 492003 329689 492037
rect 329757 492003 329769 492037
rect 329677 491997 329769 492003
rect 329804 491910 329838 492075
rect 329886 492159 329920 492334
rect 329953 492231 330045 492237
rect 329953 492197 329965 492231
rect 330033 492197 330045 492231
rect 329953 492191 330045 492197
rect 330229 492231 330321 492237
rect 330229 492197 330241 492231
rect 330309 492197 330321 492231
rect 330229 492191 330321 492197
rect 330078 492159 330108 492170
rect 329886 492147 329943 492159
rect 329886 492087 329903 492147
rect 329937 492087 329943 492147
rect 329886 492075 329943 492087
rect 330055 492147 330108 492159
rect 330055 492087 330061 492147
rect 330095 492087 330108 492147
rect 330055 492075 330108 492087
rect 329886 492072 329920 492075
rect 329953 492037 330045 492043
rect 329953 492003 329965 492037
rect 330033 492003 330045 492037
rect 329953 491997 330045 492003
rect 330078 491910 330108 492075
rect 330166 492159 330196 492172
rect 330356 492159 330390 492334
rect 330166 492147 330219 492159
rect 330166 492087 330179 492147
rect 330213 492087 330219 492147
rect 330166 492075 330219 492087
rect 330331 492147 330390 492159
rect 330331 492087 330337 492147
rect 330371 492087 330390 492147
rect 330331 492075 330390 492087
rect 330166 491910 330196 492075
rect 330356 492074 330390 492075
rect 330442 492159 330476 492334
rect 330505 492231 330597 492237
rect 330505 492197 330517 492231
rect 330585 492197 330597 492231
rect 330505 492191 330597 492197
rect 330781 492231 330873 492237
rect 330781 492197 330793 492231
rect 330861 492197 330873 492231
rect 330781 492191 330873 492197
rect 330626 492159 330656 492172
rect 330442 492147 330495 492159
rect 330442 492087 330455 492147
rect 330489 492087 330495 492147
rect 330442 492075 330495 492087
rect 330607 492147 330656 492159
rect 330607 492087 330613 492147
rect 330647 492087 330656 492147
rect 330607 492075 330656 492087
rect 330442 492068 330476 492075
rect 330229 492037 330321 492043
rect 330229 492003 330241 492037
rect 330309 492003 330321 492037
rect 330229 491997 330321 492003
rect 330505 492037 330597 492043
rect 330505 492003 330517 492037
rect 330585 492003 330597 492037
rect 330505 491997 330597 492003
rect 330626 491910 330656 492075
rect 330718 492159 330748 492172
rect 330908 492159 330942 492334
rect 330718 492147 330771 492159
rect 330718 492087 330731 492147
rect 330765 492087 330771 492147
rect 330718 492075 330771 492087
rect 330883 492147 330942 492159
rect 330883 492087 330889 492147
rect 330923 492087 330942 492147
rect 330883 492076 330942 492087
rect 330994 492159 331028 492334
rect 331057 492231 331149 492237
rect 331057 492197 331069 492231
rect 331137 492197 331149 492231
rect 331057 492191 331149 492197
rect 331333 492231 331425 492237
rect 331333 492197 331345 492231
rect 331413 492197 331425 492231
rect 331333 492191 331425 492197
rect 331180 492159 331210 492172
rect 330994 492147 331047 492159
rect 330994 492087 331007 492147
rect 331041 492087 331047 492147
rect 330883 492075 330929 492076
rect 330994 492075 331047 492087
rect 331159 492147 331210 492159
rect 331159 492087 331165 492147
rect 331199 492087 331210 492147
rect 331159 492075 331210 492087
rect 330718 491910 330748 492075
rect 330994 492072 331028 492075
rect 330781 492037 330873 492043
rect 330781 492003 330793 492037
rect 330861 492003 330873 492037
rect 330781 491997 330873 492003
rect 331057 492037 331149 492043
rect 331057 492003 331069 492037
rect 331137 492003 331149 492037
rect 331057 491997 331149 492003
rect 331180 491910 331210 492075
rect 331272 492159 331302 492172
rect 331458 492159 331492 492334
rect 331272 492147 331323 492159
rect 331272 492087 331283 492147
rect 331317 492087 331323 492147
rect 331272 492075 331323 492087
rect 331435 492147 331492 492159
rect 331435 492087 331441 492147
rect 331475 492087 331492 492147
rect 331435 492075 331492 492087
rect 331272 491910 331302 492075
rect 331458 492072 331492 492075
rect 331546 492159 331580 492334
rect 331609 492231 331701 492237
rect 331609 492197 331621 492231
rect 331689 492197 331701 492231
rect 331609 492191 331701 492197
rect 331885 492231 331977 492237
rect 331885 492197 331897 492231
rect 331965 492197 331977 492231
rect 331885 492191 331977 492197
rect 331732 492159 331762 492172
rect 331546 492147 331599 492159
rect 331546 492087 331559 492147
rect 331593 492087 331599 492147
rect 331546 492075 331599 492087
rect 331711 492147 331762 492159
rect 331711 492087 331717 492147
rect 331751 492087 331762 492147
rect 331711 492075 331762 492087
rect 331546 492070 331580 492075
rect 331333 492037 331425 492043
rect 331333 492003 331345 492037
rect 331413 492003 331425 492037
rect 331333 491997 331425 492003
rect 331609 492037 331701 492043
rect 331609 492003 331621 492037
rect 331689 492003 331701 492037
rect 331609 491997 331701 492003
rect 331732 491910 331762 492075
rect 331818 492159 331848 492172
rect 332014 492159 332048 492334
rect 331818 492147 331875 492159
rect 331818 492087 331835 492147
rect 331869 492087 331875 492147
rect 331818 492075 331875 492087
rect 331987 492147 332048 492159
rect 331987 492087 331993 492147
rect 332027 492087 332048 492147
rect 331987 492075 332048 492087
rect 331818 491910 331848 492075
rect 332014 492066 332048 492075
rect 332096 492159 332130 492334
rect 332161 492231 332253 492237
rect 332161 492197 332173 492231
rect 332241 492197 332253 492231
rect 332161 492191 332253 492197
rect 332437 492231 332529 492237
rect 332437 492197 332449 492231
rect 332517 492197 332529 492231
rect 332437 492191 332529 492197
rect 332286 492159 332316 492172
rect 332096 492147 332151 492159
rect 332096 492087 332111 492147
rect 332145 492087 332151 492147
rect 332096 492075 332151 492087
rect 332263 492147 332316 492159
rect 332263 492087 332269 492147
rect 332303 492087 332316 492147
rect 332263 492075 332316 492087
rect 332096 492072 332130 492075
rect 331885 492037 331977 492043
rect 331885 492003 331897 492037
rect 331965 492003 331977 492037
rect 331885 491997 331977 492003
rect 332161 492037 332253 492043
rect 332161 492003 332173 492037
rect 332241 492003 332253 492037
rect 332161 491997 332253 492003
rect 332286 491910 332316 492075
rect 332374 492159 332404 492170
rect 332568 492159 332602 492334
rect 332374 492147 332427 492159
rect 332374 492087 332387 492147
rect 332421 492087 332427 492147
rect 332374 492075 332427 492087
rect 332539 492147 332602 492159
rect 332539 492087 332545 492147
rect 332579 492087 332602 492147
rect 332539 492075 332602 492087
rect 332374 491910 332404 492075
rect 332568 492070 332602 492075
rect 332646 492159 332680 492334
rect 332713 492231 332805 492237
rect 332713 492197 332725 492231
rect 332793 492197 332805 492231
rect 332713 492191 332805 492197
rect 332989 492231 333081 492237
rect 332989 492197 333001 492231
rect 333069 492197 333081 492231
rect 332989 492191 333081 492197
rect 332838 492159 332868 492174
rect 332646 492147 332703 492159
rect 332646 492087 332663 492147
rect 332697 492087 332703 492147
rect 332646 492075 332703 492087
rect 332815 492147 332868 492159
rect 332815 492087 332821 492147
rect 332855 492087 332868 492147
rect 332815 492075 332868 492087
rect 332646 492072 332680 492075
rect 332437 492037 332529 492043
rect 332437 492003 332449 492037
rect 332517 492003 332529 492037
rect 332437 491997 332529 492003
rect 332713 492037 332805 492043
rect 332713 492003 332725 492037
rect 332793 492003 332805 492037
rect 332713 491997 332805 492003
rect 332838 491910 332868 492075
rect 332926 492159 332956 492174
rect 333124 492159 333158 492334
rect 332926 492147 332979 492159
rect 332926 492087 332939 492147
rect 332973 492087 332979 492147
rect 332926 492075 332979 492087
rect 333091 492147 333158 492159
rect 333091 492087 333097 492147
rect 333131 492087 333158 492147
rect 333091 492075 333158 492087
rect 332926 491910 332956 492075
rect 333124 492062 333158 492075
rect 333198 492159 333232 492334
rect 333265 492231 333357 492237
rect 333265 492197 333277 492231
rect 333345 492197 333357 492231
rect 333265 492191 333357 492197
rect 333541 492231 333633 492237
rect 333541 492197 333553 492231
rect 333621 492197 333633 492231
rect 333541 492191 333633 492197
rect 333388 492159 333418 492176
rect 333198 492147 333255 492159
rect 333198 492087 333215 492147
rect 333249 492087 333255 492147
rect 333198 492075 333255 492087
rect 333367 492147 333418 492159
rect 333367 492087 333373 492147
rect 333407 492087 333418 492147
rect 333367 492075 333418 492087
rect 333198 492066 333232 492075
rect 332989 492037 333081 492043
rect 332989 492003 333001 492037
rect 333069 492003 333081 492037
rect 332989 491997 333081 492003
rect 333265 492037 333357 492043
rect 333265 492003 333277 492037
rect 333345 492003 333357 492037
rect 333265 491997 333357 492003
rect 333388 491910 333418 492075
rect 333476 492159 333506 492174
rect 333668 492159 333702 492334
rect 333476 492147 333531 492159
rect 333476 492087 333491 492147
rect 333525 492087 333531 492147
rect 333476 492075 333531 492087
rect 333643 492147 333702 492159
rect 333643 492087 333649 492147
rect 333683 492087 333702 492147
rect 333643 492075 333702 492087
rect 333476 491910 333506 492075
rect 333668 492062 333702 492075
rect 333748 492159 333782 492334
rect 333817 492231 333909 492237
rect 333817 492197 333829 492231
rect 333897 492197 333909 492231
rect 333817 492191 333909 492197
rect 334093 492231 334185 492237
rect 334093 492197 334105 492231
rect 334173 492197 334185 492231
rect 334093 492191 334185 492197
rect 333940 492159 333970 492174
rect 333748 492147 333807 492159
rect 333748 492087 333767 492147
rect 333801 492087 333807 492147
rect 333748 492075 333807 492087
rect 333919 492147 333970 492159
rect 333919 492087 333925 492147
rect 333959 492087 333970 492147
rect 333919 492075 333970 492087
rect 333748 492060 333782 492075
rect 333541 492037 333633 492043
rect 333541 492003 333553 492037
rect 333621 492003 333633 492037
rect 333541 491997 333633 492003
rect 333817 492037 333909 492043
rect 333817 492003 333829 492037
rect 333897 492003 333909 492037
rect 333817 491997 333909 492003
rect 333940 491910 333970 492075
rect 334028 492159 334058 492176
rect 334224 492159 334258 492334
rect 334028 492147 334083 492159
rect 334028 492087 334043 492147
rect 334077 492087 334083 492147
rect 334028 492075 334083 492087
rect 334195 492147 334258 492159
rect 334195 492087 334201 492147
rect 334235 492087 334258 492147
rect 334195 492075 334258 492087
rect 334028 491910 334058 492075
rect 334224 492062 334258 492075
rect 334298 492159 334332 492334
rect 334369 492231 334461 492237
rect 334369 492197 334381 492231
rect 334449 492197 334461 492231
rect 334369 492191 334461 492197
rect 334645 492231 334737 492237
rect 334645 492197 334657 492231
rect 334725 492197 334737 492231
rect 334645 492191 334737 492197
rect 334492 492159 334522 492174
rect 334298 492147 334359 492159
rect 334298 492087 334319 492147
rect 334353 492087 334359 492147
rect 334298 492075 334359 492087
rect 334471 492147 334522 492159
rect 334471 492087 334477 492147
rect 334511 492087 334522 492147
rect 334471 492075 334522 492087
rect 334298 492060 334332 492075
rect 334093 492037 334185 492043
rect 334093 492003 334105 492037
rect 334173 492003 334185 492037
rect 334093 491997 334185 492003
rect 334369 492037 334461 492043
rect 334369 492003 334381 492037
rect 334449 492003 334461 492037
rect 334369 491997 334461 492003
rect 334492 491910 334522 492075
rect 334582 492159 334612 492176
rect 334774 492159 334808 492334
rect 334582 492147 334635 492159
rect 334582 492087 334595 492147
rect 334629 492087 334635 492147
rect 334582 492075 334635 492087
rect 334747 492147 334808 492159
rect 334747 492087 334753 492147
rect 334787 492087 334808 492147
rect 334747 492075 334808 492087
rect 334582 491910 334612 492075
rect 334774 492064 334808 492075
rect 334850 492159 334884 492334
rect 334921 492231 335013 492237
rect 334921 492197 334933 492231
rect 335001 492197 335013 492231
rect 334921 492191 335013 492197
rect 335197 492231 335289 492237
rect 335197 492197 335209 492231
rect 335277 492197 335289 492231
rect 335197 492191 335289 492197
rect 335044 492159 335074 492174
rect 334850 492147 334911 492159
rect 334850 492087 334871 492147
rect 334905 492087 334911 492147
rect 334850 492075 334911 492087
rect 335023 492147 335074 492159
rect 335023 492087 335029 492147
rect 335063 492087 335074 492147
rect 335023 492075 335074 492087
rect 334850 492064 334884 492075
rect 334645 492037 334737 492043
rect 334645 492003 334657 492037
rect 334725 492003 334737 492037
rect 334645 491997 334737 492003
rect 334921 492037 335013 492043
rect 334921 492003 334933 492037
rect 335001 492003 335013 492037
rect 334921 491997 335013 492003
rect 335044 491910 335074 492075
rect 335134 492159 335164 492176
rect 335324 492159 335358 492334
rect 335134 492147 335187 492159
rect 335134 492087 335147 492147
rect 335181 492087 335187 492147
rect 335134 492075 335187 492087
rect 335299 492147 335358 492159
rect 335299 492087 335305 492147
rect 335339 492087 335358 492147
rect 335299 492075 335358 492087
rect 335134 491910 335164 492075
rect 335324 492068 335358 492075
rect 335406 492159 335440 492334
rect 335473 492231 335565 492237
rect 335473 492197 335485 492231
rect 335553 492197 335565 492231
rect 335473 492191 335565 492197
rect 335749 492231 335841 492237
rect 335749 492197 335761 492231
rect 335829 492197 335841 492231
rect 335749 492191 335841 492197
rect 335598 492159 335628 492180
rect 335406 492147 335463 492159
rect 335406 492087 335423 492147
rect 335457 492087 335463 492147
rect 335406 492075 335463 492087
rect 335575 492147 335628 492159
rect 335575 492087 335581 492147
rect 335615 492087 335628 492147
rect 335575 492075 335628 492087
rect 335406 492066 335440 492075
rect 335197 492037 335289 492043
rect 335197 492003 335209 492037
rect 335277 492003 335289 492037
rect 335197 491997 335289 492003
rect 335473 492037 335565 492043
rect 335473 492003 335485 492037
rect 335553 492003 335565 492037
rect 335473 491997 335565 492003
rect 335598 491910 335628 492075
rect 335688 492159 335718 492182
rect 335876 492159 335910 492334
rect 335688 492147 335739 492159
rect 335688 492087 335699 492147
rect 335733 492087 335739 492147
rect 335688 492075 335739 492087
rect 335851 492147 335910 492159
rect 335851 492087 335857 492147
rect 335891 492087 335910 492147
rect 335851 492075 335910 492087
rect 335688 491910 335718 492075
rect 335876 492072 335910 492075
rect 335954 492159 335988 492334
rect 336025 492231 336117 492237
rect 336025 492197 336037 492231
rect 336105 492197 336117 492231
rect 336025 492191 336117 492197
rect 336301 492231 336393 492237
rect 336301 492197 336313 492231
rect 336381 492197 336393 492231
rect 336301 492191 336393 492197
rect 336152 492159 336182 492182
rect 335954 492147 336015 492159
rect 335954 492087 335975 492147
rect 336009 492087 336015 492147
rect 335954 492075 336015 492087
rect 336127 492147 336182 492159
rect 336127 492087 336133 492147
rect 336167 492087 336182 492147
rect 336127 492075 336182 492087
rect 335954 492074 335988 492075
rect 335749 492037 335841 492043
rect 335749 492003 335761 492037
rect 335829 492003 335841 492037
rect 335749 491997 335841 492003
rect 336025 492037 336117 492043
rect 336025 492003 336037 492037
rect 336105 492003 336117 492037
rect 336025 491997 336117 492003
rect 336152 491910 336182 492075
rect 336238 492159 336268 492186
rect 336426 492159 336460 492334
rect 336238 492147 336291 492159
rect 336238 492087 336251 492147
rect 336285 492087 336291 492147
rect 336238 492075 336291 492087
rect 336403 492147 336460 492159
rect 336403 492087 336409 492147
rect 336443 492087 336460 492147
rect 336403 492075 336460 492087
rect 336238 491910 336268 492075
rect 336426 492070 336460 492075
rect 336510 492159 336544 492334
rect 336577 492231 336669 492237
rect 336577 492197 336589 492231
rect 336657 492197 336669 492231
rect 336577 492191 336669 492197
rect 336853 492231 336945 492237
rect 336853 492197 336865 492231
rect 336933 492197 336945 492231
rect 336853 492191 336945 492197
rect 336698 492159 336728 492172
rect 336510 492147 336567 492159
rect 336510 492087 336527 492147
rect 336561 492087 336567 492147
rect 336510 492075 336567 492087
rect 336679 492147 336728 492159
rect 336679 492087 336685 492147
rect 336719 492087 336728 492147
rect 336679 492075 336728 492087
rect 336510 492068 336544 492075
rect 336301 492037 336393 492043
rect 336301 492003 336313 492037
rect 336381 492003 336393 492037
rect 336301 491997 336393 492003
rect 336577 492037 336669 492043
rect 336577 492003 336589 492037
rect 336657 492003 336669 492037
rect 336577 491997 336669 492003
rect 336698 491910 336728 492075
rect 336790 492159 336820 492170
rect 336978 492159 337012 492334
rect 336790 492147 336843 492159
rect 336790 492087 336803 492147
rect 336837 492087 336843 492147
rect 336790 492075 336843 492087
rect 336955 492147 337012 492159
rect 336955 492087 336961 492147
rect 336995 492087 337012 492147
rect 336955 492075 337012 492087
rect 336790 491910 336820 492075
rect 336978 492070 337012 492075
rect 337062 492159 337096 492334
rect 337129 492231 337221 492237
rect 337129 492197 337141 492231
rect 337209 492197 337221 492231
rect 337129 492191 337221 492197
rect 337405 492231 337497 492237
rect 337405 492197 337417 492231
rect 337485 492197 337497 492231
rect 337405 492191 337497 492197
rect 337254 492159 337284 492172
rect 337062 492147 337119 492159
rect 337062 492087 337079 492147
rect 337113 492087 337119 492147
rect 337062 492075 337119 492087
rect 337231 492147 337284 492159
rect 337231 492087 337237 492147
rect 337271 492087 337284 492147
rect 337231 492075 337284 492087
rect 337062 492072 337096 492075
rect 336853 492037 336945 492043
rect 336853 492003 336865 492037
rect 336933 492003 336945 492037
rect 336853 491997 336945 492003
rect 337129 492037 337221 492043
rect 337129 492003 337141 492037
rect 337209 492003 337221 492037
rect 337129 491997 337221 492003
rect 337254 491910 337284 492075
rect 337338 492159 337368 492172
rect 337532 492159 337566 492334
rect 337338 492147 337395 492159
rect 337338 492087 337355 492147
rect 337389 492087 337395 492147
rect 337338 492075 337395 492087
rect 337507 492147 337566 492159
rect 337507 492087 337513 492147
rect 337547 492087 337566 492147
rect 337507 492076 337566 492087
rect 337610 492159 337644 492334
rect 337681 492231 337773 492237
rect 337681 492197 337693 492231
rect 337761 492197 337773 492231
rect 337681 492191 337773 492197
rect 337804 492159 337834 492172
rect 337610 492147 337671 492159
rect 337610 492087 337631 492147
rect 337665 492087 337671 492147
rect 337507 492075 337553 492076
rect 337610 492075 337671 492087
rect 337783 492147 337834 492159
rect 337783 492087 337789 492147
rect 337823 492087 337834 492147
rect 337783 492075 337834 492087
rect 337924 492082 337958 492334
rect 337338 491910 337368 492075
rect 337610 492074 337644 492075
rect 337405 492037 337497 492043
rect 337405 492003 337417 492037
rect 337485 492003 337497 492037
rect 337405 491997 337497 492003
rect 337681 492037 337773 492043
rect 337681 492003 337693 492037
rect 337761 492003 337773 492037
rect 337681 491997 337773 492003
rect 337804 491910 337834 492075
rect 323667 491868 337836 491910
rect 337794 491866 337836 491868
rect 158318 491723 159188 491755
rect 143461 491657 159188 491723
rect 143341 491553 143433 491559
rect 143341 491519 143353 491553
rect 143421 491519 143433 491553
rect 143341 491513 143433 491519
rect 143466 491481 143506 491657
rect 143285 491469 143331 491481
rect 58039 491388 61532 491434
rect 141258 491411 143291 491469
rect 61030 491386 61062 491388
rect 59538 491334 59660 491344
rect 59538 491290 59566 491334
rect 59638 491290 59660 491334
rect 59538 491108 59660 491290
rect 60000 491270 60090 491286
rect 60000 491206 60012 491270
rect 60084 491206 60090 491270
rect 59504 491100 59704 491108
rect 58428 490908 59704 491100
rect 58428 490882 59702 490908
rect 52872 490836 59702 490882
rect 52872 490618 58692 490836
rect 52872 489146 53136 490618
rect 60000 490340 60090 491206
rect 57078 490336 59388 490340
rect 59652 490336 61758 490340
rect 57078 489740 61758 490336
rect 52310 480230 53762 489146
rect 57078 488820 58038 489740
rect 57078 488220 57238 488820
rect 57838 488220 58038 488820
rect 57078 488060 58038 488220
rect 60798 488820 61758 489740
rect 60798 488220 60958 488820
rect 61558 488220 61758 488820
rect 141258 489730 142348 491411
rect 143127 491233 143169 491411
rect 143285 491409 143291 491411
rect 143325 491409 143331 491469
rect 143285 491397 143331 491409
rect 143443 491469 143506 491481
rect 143443 491409 143449 491469
rect 143483 491409 143506 491469
rect 143443 491397 143506 491409
rect 143466 491391 143506 491397
rect 143548 491481 143588 491657
rect 143617 491553 143709 491559
rect 143617 491519 143629 491553
rect 143697 491519 143709 491553
rect 143617 491513 143709 491519
rect 143893 491553 143985 491559
rect 143893 491519 143905 491553
rect 143973 491519 143985 491553
rect 143893 491513 143985 491519
rect 143742 491481 143772 491489
rect 143548 491469 143607 491481
rect 143548 491409 143567 491469
rect 143601 491409 143607 491469
rect 143548 491397 143607 491409
rect 143719 491469 143772 491481
rect 143719 491409 143725 491469
rect 143759 491409 143772 491469
rect 143719 491397 143772 491409
rect 143548 491393 143588 491397
rect 143341 491359 143433 491365
rect 143341 491325 143353 491359
rect 143421 491325 143433 491359
rect 143341 491319 143433 491325
rect 143617 491359 143709 491365
rect 143617 491325 143629 491359
rect 143697 491325 143709 491359
rect 143617 491319 143709 491325
rect 143742 491233 143772 491397
rect 143828 491481 143858 491489
rect 144024 491481 144064 491657
rect 143828 491469 143883 491481
rect 143828 491409 143843 491469
rect 143877 491409 143883 491469
rect 143828 491397 143883 491409
rect 143995 491469 144064 491481
rect 143995 491409 144001 491469
rect 144035 491409 144064 491469
rect 143995 491397 144064 491409
rect 143828 491233 143858 491397
rect 144024 491393 144064 491397
rect 144092 491481 144132 491657
rect 144169 491553 144261 491559
rect 144169 491519 144181 491553
rect 144249 491519 144261 491553
rect 144169 491513 144261 491519
rect 144445 491553 144537 491559
rect 144445 491519 144457 491553
rect 144525 491519 144537 491553
rect 144445 491513 144537 491519
rect 144296 491481 144326 491489
rect 144092 491469 144159 491481
rect 144092 491409 144119 491469
rect 144153 491409 144159 491469
rect 144092 491397 144159 491409
rect 144271 491469 144326 491481
rect 144271 491409 144277 491469
rect 144311 491409 144326 491469
rect 144271 491397 144326 491409
rect 144092 491393 144132 491397
rect 143893 491359 143985 491365
rect 143893 491325 143905 491359
rect 143973 491325 143985 491359
rect 143893 491319 143985 491325
rect 144169 491359 144261 491365
rect 144169 491325 144181 491359
rect 144249 491325 144261 491359
rect 144169 491319 144261 491325
rect 144296 491233 144326 491397
rect 144382 491481 144412 491489
rect 144572 491481 144612 491657
rect 144382 491469 144435 491481
rect 144382 491409 144395 491469
rect 144429 491409 144435 491469
rect 144382 491397 144435 491409
rect 144547 491469 144612 491481
rect 144547 491409 144553 491469
rect 144587 491409 144612 491469
rect 144547 491397 144612 491409
rect 144382 491233 144412 491397
rect 144572 491389 144612 491397
rect 144644 491481 144684 491657
rect 144721 491553 144813 491559
rect 144721 491519 144733 491553
rect 144801 491519 144813 491553
rect 144721 491513 144813 491519
rect 144997 491553 145089 491559
rect 144997 491519 145009 491553
rect 145077 491519 145089 491553
rect 144997 491513 145089 491519
rect 144844 491481 144874 491489
rect 144644 491469 144711 491481
rect 144644 491409 144671 491469
rect 144705 491409 144711 491469
rect 144644 491397 144711 491409
rect 144823 491469 144874 491481
rect 144823 491409 144829 491469
rect 144863 491409 144874 491469
rect 144823 491397 144874 491409
rect 144644 491393 144684 491397
rect 144445 491359 144537 491365
rect 144445 491325 144457 491359
rect 144525 491325 144537 491359
rect 144445 491319 144537 491325
rect 144721 491359 144813 491365
rect 144721 491325 144733 491359
rect 144801 491325 144813 491359
rect 144721 491319 144813 491325
rect 144844 491233 144874 491397
rect 144936 491481 144966 491487
rect 145124 491481 145164 491657
rect 144936 491469 144987 491481
rect 144936 491409 144947 491469
rect 144981 491409 144987 491469
rect 144936 491397 144987 491409
rect 145099 491469 145164 491481
rect 145099 491409 145105 491469
rect 145139 491409 145164 491469
rect 145099 491397 145164 491409
rect 145204 491481 145244 491657
rect 145273 491553 145365 491559
rect 145273 491519 145285 491553
rect 145353 491519 145365 491553
rect 145273 491513 145365 491519
rect 145549 491553 145641 491559
rect 145549 491519 145561 491553
rect 145629 491519 145641 491553
rect 145549 491513 145641 491519
rect 145394 491481 145424 491487
rect 145204 491469 145263 491481
rect 145204 491409 145223 491469
rect 145257 491409 145263 491469
rect 145204 491397 145263 491409
rect 145375 491469 145424 491481
rect 145375 491409 145381 491469
rect 145415 491409 145424 491469
rect 145375 491397 145424 491409
rect 144936 491233 144966 491397
rect 144997 491359 145089 491365
rect 144997 491325 145009 491359
rect 145077 491325 145089 491359
rect 144997 491319 145089 491325
rect 145273 491359 145365 491365
rect 145273 491325 145285 491359
rect 145353 491325 145365 491359
rect 145273 491319 145365 491325
rect 145394 491233 145424 491397
rect 145486 491481 145516 491485
rect 145678 491481 145718 491657
rect 145486 491469 145539 491481
rect 145486 491409 145499 491469
rect 145533 491409 145539 491469
rect 145486 491397 145539 491409
rect 145651 491469 145718 491481
rect 145651 491409 145657 491469
rect 145691 491409 145718 491469
rect 145651 491397 145718 491409
rect 145486 491233 145516 491397
rect 145678 491393 145718 491397
rect 145752 491481 145792 491657
rect 145825 491553 145917 491559
rect 145825 491519 145837 491553
rect 145905 491519 145917 491553
rect 145825 491513 145917 491519
rect 146101 491553 146193 491559
rect 146101 491519 146113 491553
rect 146181 491519 146193 491553
rect 146101 491513 146193 491519
rect 145950 491481 145980 491485
rect 145752 491469 145815 491481
rect 145752 491409 145775 491469
rect 145809 491409 145815 491469
rect 145752 491397 145815 491409
rect 145927 491469 145980 491481
rect 145927 491409 145933 491469
rect 145967 491409 145980 491469
rect 145927 491397 145980 491409
rect 145752 491395 145792 491397
rect 145549 491359 145641 491365
rect 145549 491325 145561 491359
rect 145629 491325 145641 491359
rect 145549 491319 145641 491325
rect 145825 491359 145917 491365
rect 145825 491325 145837 491359
rect 145905 491325 145917 491359
rect 145825 491319 145917 491325
rect 145950 491233 145980 491397
rect 146038 491481 146068 491483
rect 146230 491481 146270 491657
rect 146038 491469 146091 491481
rect 146038 491409 146051 491469
rect 146085 491409 146091 491469
rect 146038 491397 146091 491409
rect 146203 491469 146270 491481
rect 146203 491409 146209 491469
rect 146243 491409 146270 491469
rect 146203 491397 146270 491409
rect 146038 491233 146068 491397
rect 146230 491391 146270 491397
rect 146300 491481 146340 491657
rect 146377 491553 146469 491559
rect 146377 491519 146389 491553
rect 146457 491519 146469 491553
rect 146377 491513 146469 491519
rect 146653 491553 146745 491559
rect 146653 491519 146665 491553
rect 146733 491519 146745 491553
rect 146653 491513 146745 491519
rect 146500 491481 146530 491483
rect 146300 491469 146367 491481
rect 146300 491409 146327 491469
rect 146361 491409 146367 491469
rect 146300 491397 146367 491409
rect 146479 491469 146530 491481
rect 146479 491409 146485 491469
rect 146519 491409 146530 491469
rect 146479 491397 146530 491409
rect 146300 491395 146340 491397
rect 146101 491359 146193 491365
rect 146377 491363 146469 491365
rect 146101 491325 146113 491359
rect 146181 491325 146193 491359
rect 146374 491359 146469 491363
rect 146374 491330 146389 491359
rect 146101 491319 146193 491325
rect 146377 491325 146389 491330
rect 146457 491325 146469 491359
rect 146377 491319 146469 491325
rect 146500 491233 146530 491397
rect 146588 491481 146618 491483
rect 146778 491481 146818 491657
rect 146588 491469 146643 491481
rect 146588 491409 146603 491469
rect 146637 491409 146643 491469
rect 146588 491397 146643 491409
rect 146755 491469 146818 491481
rect 146755 491409 146761 491469
rect 146795 491409 146818 491469
rect 146755 491397 146818 491409
rect 146588 491233 146618 491397
rect 146778 491391 146818 491397
rect 146856 491481 146896 491657
rect 146929 491553 147021 491559
rect 146929 491519 146941 491553
rect 147009 491519 147021 491553
rect 146929 491513 147021 491519
rect 147205 491553 147297 491559
rect 147205 491519 147217 491553
rect 147285 491519 147297 491553
rect 147205 491513 147297 491519
rect 147052 491481 147082 491485
rect 146856 491469 146919 491481
rect 146856 491409 146879 491469
rect 146913 491409 146919 491469
rect 146856 491397 146919 491409
rect 147031 491469 147082 491481
rect 147031 491409 147037 491469
rect 147071 491409 147082 491469
rect 147031 491397 147082 491409
rect 146856 491395 146896 491397
rect 146653 491359 146745 491365
rect 146653 491325 146665 491359
rect 146733 491325 146745 491359
rect 146653 491319 146745 491325
rect 146929 491359 147021 491365
rect 146929 491325 146941 491359
rect 147009 491325 147021 491359
rect 146929 491319 147021 491325
rect 147052 491233 147082 491397
rect 147140 491481 147170 491485
rect 147332 491481 147372 491657
rect 147140 491469 147195 491481
rect 147140 491409 147155 491469
rect 147189 491409 147195 491469
rect 147140 491397 147195 491409
rect 147307 491469 147372 491481
rect 147307 491409 147313 491469
rect 147347 491409 147372 491469
rect 147307 491397 147372 491409
rect 147140 491233 147170 491397
rect 147332 491383 147372 491397
rect 147410 491481 147450 491657
rect 147481 491553 147573 491559
rect 147481 491519 147493 491553
rect 147561 491519 147573 491553
rect 147481 491513 147573 491519
rect 147757 491553 147849 491559
rect 147757 491519 147769 491553
rect 147837 491519 147849 491553
rect 147757 491513 147849 491519
rect 147604 491481 147634 491485
rect 147410 491469 147471 491481
rect 147410 491409 147431 491469
rect 147465 491409 147471 491469
rect 147410 491397 147471 491409
rect 147583 491469 147634 491481
rect 147583 491409 147589 491469
rect 147623 491409 147634 491469
rect 147583 491397 147634 491409
rect 147410 491391 147450 491397
rect 147205 491359 147297 491365
rect 147205 491325 147217 491359
rect 147285 491325 147297 491359
rect 147205 491319 147297 491325
rect 147481 491359 147573 491365
rect 147481 491325 147493 491359
rect 147561 491325 147573 491359
rect 147481 491319 147573 491325
rect 147604 491233 147634 491397
rect 147696 491481 147726 491485
rect 147888 491481 147928 491657
rect 147696 491469 147747 491481
rect 147696 491409 147707 491469
rect 147741 491409 147747 491469
rect 147696 491397 147747 491409
rect 147859 491469 147928 491481
rect 147859 491409 147865 491469
rect 147899 491409 147928 491469
rect 147859 491397 147928 491409
rect 147962 491481 148002 491657
rect 148033 491553 148125 491559
rect 148033 491519 148045 491553
rect 148113 491519 148125 491553
rect 148033 491513 148125 491519
rect 148309 491553 148401 491559
rect 148309 491519 148321 491553
rect 148389 491519 148401 491553
rect 148309 491513 148401 491519
rect 148158 491481 148188 491495
rect 147962 491469 148023 491481
rect 147962 491409 147983 491469
rect 148017 491409 148023 491469
rect 147962 491397 148023 491409
rect 148135 491469 148188 491481
rect 148135 491409 148141 491469
rect 148175 491409 148188 491469
rect 148135 491397 148188 491409
rect 147696 491233 147726 491397
rect 147888 491393 147928 491397
rect 147757 491359 147849 491365
rect 147757 491325 147769 491359
rect 147837 491325 147849 491359
rect 147757 491319 147849 491325
rect 148033 491359 148125 491365
rect 148033 491325 148045 491359
rect 148113 491325 148125 491359
rect 148033 491319 148125 491325
rect 148158 491233 148188 491397
rect 148244 491481 148274 491493
rect 148432 491481 148466 491657
rect 148244 491469 148299 491481
rect 148244 491409 148259 491469
rect 148293 491409 148299 491469
rect 148244 491397 148299 491409
rect 148411 491469 148466 491481
rect 148411 491409 148417 491469
rect 148451 491409 148466 491469
rect 148411 491397 148466 491409
rect 148244 491233 148274 491397
rect 148432 491393 148466 491397
rect 148522 491481 148556 491657
rect 148585 491553 148677 491559
rect 148585 491519 148597 491553
rect 148665 491519 148677 491553
rect 148585 491513 148677 491519
rect 148861 491553 148953 491559
rect 148861 491519 148873 491553
rect 148941 491519 148953 491553
rect 148861 491513 148953 491519
rect 148712 491481 148742 491491
rect 148522 491469 148575 491481
rect 148522 491409 148535 491469
rect 148569 491409 148575 491469
rect 148522 491397 148575 491409
rect 148687 491469 148742 491481
rect 148687 491409 148693 491469
rect 148727 491409 148742 491469
rect 148687 491397 148742 491409
rect 148522 491393 148556 491397
rect 148309 491359 148401 491365
rect 148309 491325 148321 491359
rect 148389 491325 148401 491359
rect 148309 491319 148401 491325
rect 148585 491359 148677 491365
rect 148585 491325 148597 491359
rect 148665 491325 148677 491359
rect 148585 491319 148677 491325
rect 148712 491233 148742 491397
rect 148798 491481 148828 491491
rect 148988 491481 149022 491657
rect 148798 491469 148851 491481
rect 148798 491409 148811 491469
rect 148845 491409 148851 491469
rect 148798 491397 148851 491409
rect 148963 491469 149022 491481
rect 148963 491409 148969 491469
rect 149003 491409 149022 491469
rect 148963 491397 149022 491409
rect 149072 491481 149106 491657
rect 149137 491553 149229 491559
rect 149137 491519 149149 491553
rect 149217 491519 149229 491553
rect 149137 491513 149229 491519
rect 149264 491481 149298 491495
rect 149072 491469 149127 491481
rect 149072 491409 149087 491469
rect 149121 491409 149127 491469
rect 149072 491397 149127 491409
rect 149239 491469 149298 491481
rect 149239 491409 149245 491469
rect 149279 491409 149298 491469
rect 149239 491397 149298 491409
rect 148798 491233 148828 491397
rect 148988 491393 149022 491397
rect 148861 491359 148953 491365
rect 148861 491325 148873 491359
rect 148941 491325 148953 491359
rect 148861 491319 148953 491325
rect 149137 491359 149229 491365
rect 149137 491325 149149 491359
rect 149217 491325 149229 491359
rect 149137 491319 149229 491325
rect 149264 491233 149298 491397
rect 149346 491481 149380 491657
rect 149413 491553 149505 491559
rect 149413 491519 149425 491553
rect 149493 491519 149505 491553
rect 149413 491513 149505 491519
rect 149689 491553 149781 491559
rect 149689 491519 149701 491553
rect 149769 491519 149781 491553
rect 149689 491513 149781 491519
rect 149538 491481 149568 491493
rect 149346 491469 149403 491481
rect 149346 491409 149363 491469
rect 149397 491409 149403 491469
rect 149346 491397 149403 491409
rect 149515 491469 149568 491481
rect 149515 491409 149521 491469
rect 149555 491409 149568 491469
rect 149515 491397 149568 491409
rect 149346 491395 149380 491397
rect 149413 491359 149505 491365
rect 149413 491325 149425 491359
rect 149493 491325 149505 491359
rect 149413 491319 149505 491325
rect 149538 491233 149568 491397
rect 149626 491481 149656 491495
rect 149816 491481 149850 491657
rect 149626 491469 149679 491481
rect 149626 491409 149639 491469
rect 149673 491409 149679 491469
rect 149626 491397 149679 491409
rect 149791 491469 149850 491481
rect 149791 491409 149797 491469
rect 149831 491409 149850 491469
rect 149791 491397 149850 491409
rect 149902 491481 149936 491657
rect 149974 491595 150189 491605
rect 149974 491559 150104 491595
rect 149965 491553 150104 491559
rect 149965 491519 149977 491553
rect 150045 491535 150104 491553
rect 150164 491535 150189 491595
rect 150045 491525 150189 491535
rect 150241 491553 150333 491559
rect 150045 491519 150057 491525
rect 149965 491513 150057 491519
rect 150241 491519 150253 491553
rect 150321 491519 150333 491553
rect 150241 491513 150333 491519
rect 150086 491481 150116 491495
rect 149902 491469 149955 491481
rect 149902 491409 149915 491469
rect 149949 491409 149955 491469
rect 149902 491397 149955 491409
rect 150067 491469 150116 491481
rect 150067 491409 150073 491469
rect 150107 491409 150116 491469
rect 150067 491397 150116 491409
rect 149626 491233 149656 491397
rect 149902 491391 149936 491397
rect 149689 491359 149781 491365
rect 149689 491325 149701 491359
rect 149769 491325 149781 491359
rect 149965 491359 150057 491365
rect 149965 491340 149977 491359
rect 149689 491319 149781 491325
rect 149829 491335 149977 491340
rect 149829 491280 149839 491335
rect 149904 491325 149977 491335
rect 150045 491325 150057 491359
rect 149904 491319 150057 491325
rect 149904 491290 150044 491319
rect 149904 491280 149914 491290
rect 149829 491275 149914 491280
rect 150086 491233 150116 491397
rect 150178 491481 150208 491495
rect 150368 491481 150402 491657
rect 150178 491469 150231 491481
rect 150178 491409 150191 491469
rect 150225 491409 150231 491469
rect 150178 491397 150231 491409
rect 150343 491469 150402 491481
rect 150343 491409 150349 491469
rect 150383 491409 150402 491469
rect 150343 491399 150402 491409
rect 150454 491481 150488 491657
rect 150517 491553 150609 491559
rect 150517 491519 150529 491553
rect 150597 491519 150609 491553
rect 150517 491513 150609 491519
rect 150793 491553 150885 491559
rect 150793 491519 150805 491553
rect 150873 491519 150885 491553
rect 150793 491513 150885 491519
rect 150640 491481 150670 491495
rect 150454 491469 150507 491481
rect 150454 491409 150467 491469
rect 150501 491409 150507 491469
rect 150343 491397 150389 491399
rect 150454 491397 150507 491409
rect 150619 491469 150670 491481
rect 150619 491409 150625 491469
rect 150659 491409 150670 491469
rect 150619 491397 150670 491409
rect 150178 491233 150208 491397
rect 150454 491395 150488 491397
rect 150241 491359 150333 491365
rect 150241 491325 150253 491359
rect 150321 491325 150333 491359
rect 150241 491319 150333 491325
rect 150517 491359 150609 491365
rect 150517 491325 150529 491359
rect 150597 491325 150609 491359
rect 150517 491319 150609 491325
rect 150640 491233 150670 491397
rect 150732 491481 150762 491495
rect 150918 491481 150952 491657
rect 150732 491469 150783 491481
rect 150732 491409 150743 491469
rect 150777 491409 150783 491469
rect 150732 491397 150783 491409
rect 150895 491469 150952 491481
rect 150895 491409 150901 491469
rect 150935 491409 150952 491469
rect 150895 491397 150952 491409
rect 150732 491233 150762 491397
rect 150918 491395 150952 491397
rect 151006 491481 151040 491657
rect 151069 491553 151161 491559
rect 151069 491519 151081 491553
rect 151149 491519 151161 491553
rect 151069 491513 151161 491519
rect 151345 491553 151437 491559
rect 151345 491519 151357 491553
rect 151425 491519 151437 491553
rect 151345 491513 151437 491519
rect 151192 491481 151222 491495
rect 151006 491469 151059 491481
rect 151006 491409 151019 491469
rect 151053 491409 151059 491469
rect 151006 491397 151059 491409
rect 151171 491469 151222 491481
rect 151171 491409 151177 491469
rect 151211 491409 151222 491469
rect 151171 491397 151222 491409
rect 151006 491393 151040 491397
rect 150793 491359 150885 491365
rect 150793 491325 150805 491359
rect 150873 491325 150885 491359
rect 150793 491319 150885 491325
rect 151069 491359 151161 491365
rect 151069 491325 151081 491359
rect 151149 491325 151161 491359
rect 151069 491319 151161 491325
rect 151192 491233 151222 491397
rect 151278 491481 151308 491495
rect 151474 491481 151508 491657
rect 151278 491469 151335 491481
rect 151278 491409 151295 491469
rect 151329 491409 151335 491469
rect 151278 491397 151335 491409
rect 151447 491469 151508 491481
rect 151447 491409 151453 491469
rect 151487 491409 151508 491469
rect 151447 491397 151508 491409
rect 151278 491233 151308 491397
rect 151474 491389 151508 491397
rect 151556 491481 151590 491657
rect 151621 491553 151713 491559
rect 151621 491519 151633 491553
rect 151701 491519 151713 491553
rect 151621 491513 151713 491519
rect 151897 491553 151989 491559
rect 151897 491519 151909 491553
rect 151977 491519 151989 491553
rect 151897 491513 151989 491519
rect 151746 491481 151776 491495
rect 151556 491469 151611 491481
rect 151556 491409 151571 491469
rect 151605 491409 151611 491469
rect 151556 491397 151611 491409
rect 151723 491469 151776 491481
rect 151723 491409 151729 491469
rect 151763 491409 151776 491469
rect 151723 491397 151776 491409
rect 151556 491395 151590 491397
rect 151345 491359 151437 491365
rect 151345 491325 151357 491359
rect 151425 491325 151437 491359
rect 151345 491319 151437 491325
rect 151621 491359 151713 491365
rect 151621 491325 151633 491359
rect 151701 491325 151713 491359
rect 151621 491319 151713 491325
rect 151746 491233 151776 491397
rect 151834 491481 151864 491493
rect 152028 491481 152062 491657
rect 151834 491469 151887 491481
rect 151834 491409 151847 491469
rect 151881 491409 151887 491469
rect 151834 491397 151887 491409
rect 151999 491469 152062 491481
rect 151999 491409 152005 491469
rect 152039 491409 152062 491469
rect 151999 491397 152062 491409
rect 151834 491233 151864 491397
rect 152028 491393 152062 491397
rect 152106 491481 152140 491657
rect 152173 491553 152265 491559
rect 152173 491519 152185 491553
rect 152253 491519 152265 491553
rect 152173 491513 152265 491519
rect 152449 491553 152541 491559
rect 152449 491519 152461 491553
rect 152529 491519 152541 491553
rect 152449 491513 152541 491519
rect 152298 491481 152328 491497
rect 152106 491469 152163 491481
rect 152106 491409 152123 491469
rect 152157 491409 152163 491469
rect 152106 491397 152163 491409
rect 152275 491469 152328 491481
rect 152275 491409 152281 491469
rect 152315 491409 152328 491469
rect 152275 491397 152328 491409
rect 152106 491395 152140 491397
rect 151897 491359 151989 491365
rect 151897 491325 151909 491359
rect 151977 491325 151989 491359
rect 151897 491319 151989 491325
rect 152173 491359 152265 491365
rect 152173 491325 152185 491359
rect 152253 491325 152265 491359
rect 152173 491319 152265 491325
rect 152298 491233 152328 491397
rect 152386 491481 152416 491497
rect 152584 491481 152618 491657
rect 152386 491469 152439 491481
rect 152386 491409 152399 491469
rect 152433 491409 152439 491469
rect 152386 491397 152439 491409
rect 152551 491469 152618 491481
rect 152551 491409 152557 491469
rect 152591 491409 152618 491469
rect 152551 491397 152618 491409
rect 152386 491233 152416 491397
rect 152584 491385 152618 491397
rect 152658 491481 152692 491657
rect 152725 491553 152817 491559
rect 152725 491519 152737 491553
rect 152805 491519 152817 491553
rect 152725 491513 152817 491519
rect 153001 491553 153093 491559
rect 153001 491519 153013 491553
rect 153081 491519 153093 491553
rect 153001 491513 153093 491519
rect 152848 491481 152878 491499
rect 152658 491469 152715 491481
rect 152658 491409 152675 491469
rect 152709 491409 152715 491469
rect 152658 491397 152715 491409
rect 152827 491469 152878 491481
rect 152827 491409 152833 491469
rect 152867 491409 152878 491469
rect 152827 491397 152878 491409
rect 152658 491389 152692 491397
rect 152449 491359 152541 491365
rect 152449 491325 152461 491359
rect 152529 491325 152541 491359
rect 152449 491319 152541 491325
rect 152725 491359 152817 491365
rect 152725 491325 152737 491359
rect 152805 491325 152817 491359
rect 152725 491319 152817 491325
rect 152848 491233 152878 491397
rect 152936 491481 152966 491497
rect 153128 491481 153162 491657
rect 152936 491469 152991 491481
rect 152936 491409 152951 491469
rect 152985 491409 152991 491469
rect 152936 491397 152991 491409
rect 153103 491469 153162 491481
rect 153103 491409 153109 491469
rect 153143 491409 153162 491469
rect 153103 491397 153162 491409
rect 152936 491233 152966 491397
rect 153128 491385 153162 491397
rect 153208 491481 153242 491657
rect 153277 491553 153369 491559
rect 153277 491519 153289 491553
rect 153357 491519 153369 491553
rect 153277 491513 153369 491519
rect 153553 491553 153645 491559
rect 153553 491519 153565 491553
rect 153633 491519 153645 491553
rect 153553 491513 153645 491519
rect 153400 491481 153430 491497
rect 153208 491469 153267 491481
rect 153208 491409 153227 491469
rect 153261 491409 153267 491469
rect 153208 491397 153267 491409
rect 153379 491469 153430 491481
rect 153379 491409 153385 491469
rect 153419 491409 153430 491469
rect 153379 491397 153430 491409
rect 153208 491383 153242 491397
rect 153001 491359 153093 491365
rect 153001 491325 153013 491359
rect 153081 491325 153093 491359
rect 153001 491319 153093 491325
rect 153277 491359 153369 491365
rect 153277 491325 153289 491359
rect 153357 491325 153369 491359
rect 153277 491319 153369 491325
rect 153400 491233 153430 491397
rect 153488 491481 153518 491499
rect 153684 491481 153718 491657
rect 153488 491469 153543 491481
rect 153488 491409 153503 491469
rect 153537 491409 153543 491469
rect 153488 491397 153543 491409
rect 153655 491469 153718 491481
rect 153655 491409 153661 491469
rect 153695 491409 153718 491469
rect 153655 491397 153718 491409
rect 153488 491233 153518 491397
rect 153684 491385 153718 491397
rect 153758 491481 153792 491657
rect 153829 491553 153921 491559
rect 153829 491519 153841 491553
rect 153909 491519 153921 491553
rect 153829 491513 153921 491519
rect 154105 491553 154197 491559
rect 154105 491519 154117 491553
rect 154185 491519 154197 491553
rect 154105 491513 154197 491519
rect 153952 491481 153982 491497
rect 153758 491469 153819 491481
rect 153758 491409 153779 491469
rect 153813 491409 153819 491469
rect 153758 491397 153819 491409
rect 153931 491469 153982 491481
rect 153931 491409 153937 491469
rect 153971 491409 153982 491469
rect 153931 491397 153982 491409
rect 153758 491383 153792 491397
rect 153553 491359 153645 491365
rect 153553 491325 153565 491359
rect 153633 491325 153645 491359
rect 153553 491319 153645 491325
rect 153829 491359 153921 491365
rect 153829 491325 153841 491359
rect 153909 491325 153921 491359
rect 153829 491319 153921 491325
rect 153952 491233 153982 491397
rect 154042 491481 154072 491499
rect 154234 491481 154268 491657
rect 154042 491469 154095 491481
rect 154042 491409 154055 491469
rect 154089 491409 154095 491469
rect 154042 491397 154095 491409
rect 154207 491469 154268 491481
rect 154207 491409 154213 491469
rect 154247 491409 154268 491469
rect 154207 491397 154268 491409
rect 154042 491233 154072 491397
rect 154234 491387 154268 491397
rect 154310 491481 154344 491657
rect 154381 491553 154473 491559
rect 154381 491519 154393 491553
rect 154461 491519 154473 491553
rect 154381 491513 154473 491519
rect 154657 491553 154749 491559
rect 154657 491519 154669 491553
rect 154737 491519 154749 491553
rect 154657 491513 154749 491519
rect 154504 491481 154534 491497
rect 154310 491469 154371 491481
rect 154310 491409 154331 491469
rect 154365 491409 154371 491469
rect 154310 491397 154371 491409
rect 154483 491469 154534 491481
rect 154483 491409 154489 491469
rect 154523 491409 154534 491469
rect 154483 491397 154534 491409
rect 154310 491387 154344 491397
rect 154105 491359 154197 491365
rect 154105 491325 154117 491359
rect 154185 491325 154197 491359
rect 154105 491319 154197 491325
rect 154381 491359 154473 491365
rect 154381 491325 154393 491359
rect 154461 491325 154473 491359
rect 154381 491319 154473 491325
rect 154504 491233 154534 491397
rect 154594 491481 154624 491499
rect 154784 491481 154818 491657
rect 154594 491469 154647 491481
rect 154594 491409 154607 491469
rect 154641 491409 154647 491469
rect 154594 491397 154647 491409
rect 154759 491469 154818 491481
rect 154759 491409 154765 491469
rect 154799 491409 154818 491469
rect 154759 491397 154818 491409
rect 154594 491233 154624 491397
rect 154784 491391 154818 491397
rect 154866 491481 154900 491657
rect 154933 491553 155025 491559
rect 154933 491519 154945 491553
rect 155013 491519 155025 491553
rect 154933 491513 155025 491519
rect 155209 491553 155301 491559
rect 155209 491519 155221 491553
rect 155289 491519 155301 491553
rect 155209 491513 155301 491519
rect 155058 491481 155088 491503
rect 154866 491469 154923 491481
rect 154866 491409 154883 491469
rect 154917 491409 154923 491469
rect 154866 491397 154923 491409
rect 155035 491469 155088 491481
rect 155035 491409 155041 491469
rect 155075 491409 155088 491469
rect 155035 491397 155088 491409
rect 154866 491389 154900 491397
rect 154657 491359 154749 491365
rect 154657 491325 154669 491359
rect 154737 491325 154749 491359
rect 154657 491319 154749 491325
rect 154933 491359 155025 491365
rect 154933 491325 154945 491359
rect 155013 491325 155025 491359
rect 154933 491319 155025 491325
rect 155058 491233 155088 491397
rect 155148 491481 155178 491505
rect 155336 491481 155370 491657
rect 155148 491469 155199 491481
rect 155148 491409 155159 491469
rect 155193 491409 155199 491469
rect 155148 491397 155199 491409
rect 155311 491469 155370 491481
rect 155311 491409 155317 491469
rect 155351 491409 155370 491469
rect 155311 491397 155370 491409
rect 155414 491481 155448 491657
rect 155485 491553 155577 491559
rect 155485 491519 155497 491553
rect 155565 491519 155577 491553
rect 155485 491513 155577 491519
rect 155761 491553 155853 491559
rect 155761 491519 155773 491553
rect 155841 491519 155853 491553
rect 155761 491513 155853 491519
rect 155612 491481 155642 491505
rect 155414 491469 155475 491481
rect 155414 491409 155435 491469
rect 155469 491409 155475 491469
rect 155414 491397 155475 491409
rect 155587 491469 155642 491481
rect 155587 491409 155593 491469
rect 155627 491409 155642 491469
rect 155587 491397 155642 491409
rect 155148 491233 155178 491397
rect 155336 491395 155370 491397
rect 155209 491359 155301 491365
rect 155209 491325 155221 491359
rect 155289 491325 155301 491359
rect 155209 491319 155301 491325
rect 155485 491359 155577 491365
rect 155485 491325 155497 491359
rect 155565 491325 155577 491359
rect 155485 491319 155577 491325
rect 155612 491233 155642 491397
rect 155698 491481 155728 491509
rect 155886 491481 155920 491657
rect 155698 491469 155751 491481
rect 155698 491409 155711 491469
rect 155745 491409 155751 491469
rect 155698 491397 155751 491409
rect 155863 491469 155920 491481
rect 155863 491409 155869 491469
rect 155903 491409 155920 491469
rect 155863 491397 155920 491409
rect 155698 491233 155728 491397
rect 155886 491393 155920 491397
rect 155970 491481 156004 491657
rect 156037 491553 156129 491559
rect 156037 491519 156049 491553
rect 156117 491519 156129 491553
rect 156037 491513 156129 491519
rect 156313 491553 156405 491559
rect 156313 491519 156325 491553
rect 156393 491519 156405 491553
rect 156313 491513 156405 491519
rect 156158 491481 156188 491495
rect 155970 491469 156027 491481
rect 155970 491409 155987 491469
rect 156021 491409 156027 491469
rect 155970 491397 156027 491409
rect 156139 491469 156188 491481
rect 156139 491409 156145 491469
rect 156179 491409 156188 491469
rect 156139 491397 156188 491409
rect 155970 491391 156004 491397
rect 155761 491359 155853 491365
rect 155761 491325 155773 491359
rect 155841 491325 155853 491359
rect 155761 491319 155853 491325
rect 156037 491359 156129 491365
rect 156037 491325 156049 491359
rect 156117 491325 156129 491359
rect 156037 491319 156129 491325
rect 156158 491233 156188 491397
rect 156250 491481 156280 491493
rect 156438 491481 156472 491657
rect 156250 491469 156303 491481
rect 156250 491409 156263 491469
rect 156297 491409 156303 491469
rect 156250 491397 156303 491409
rect 156415 491469 156472 491481
rect 156415 491409 156421 491469
rect 156455 491409 156472 491469
rect 156415 491397 156472 491409
rect 156250 491233 156280 491397
rect 156438 491393 156472 491397
rect 156522 491481 156556 491657
rect 156589 491553 156681 491559
rect 156589 491519 156601 491553
rect 156669 491519 156681 491553
rect 156589 491513 156681 491519
rect 156865 491553 156957 491559
rect 156865 491519 156877 491553
rect 156945 491519 156957 491553
rect 156865 491513 156957 491519
rect 156714 491481 156744 491495
rect 156522 491469 156579 491481
rect 156522 491409 156539 491469
rect 156573 491409 156579 491469
rect 156522 491397 156579 491409
rect 156691 491469 156744 491481
rect 156691 491409 156697 491469
rect 156731 491409 156744 491469
rect 156691 491397 156744 491409
rect 156522 491395 156556 491397
rect 156313 491359 156405 491365
rect 156313 491325 156325 491359
rect 156393 491325 156405 491359
rect 156313 491319 156405 491325
rect 156589 491359 156681 491365
rect 156589 491325 156601 491359
rect 156669 491325 156681 491359
rect 156589 491319 156681 491325
rect 156714 491233 156744 491397
rect 156798 491481 156828 491495
rect 156992 491481 157026 491657
rect 156798 491469 156855 491481
rect 156798 491409 156815 491469
rect 156849 491409 156855 491469
rect 156798 491397 156855 491409
rect 156967 491469 157026 491481
rect 156967 491409 156973 491469
rect 157007 491409 157026 491469
rect 156967 491399 157026 491409
rect 157070 491481 157104 491657
rect 157141 491553 157233 491559
rect 157141 491519 157153 491553
rect 157221 491519 157233 491553
rect 157141 491513 157233 491519
rect 157264 491481 157294 491495
rect 157070 491469 157131 491481
rect 157070 491409 157091 491469
rect 157125 491409 157131 491469
rect 156967 491397 157013 491399
rect 157070 491397 157131 491409
rect 157243 491469 157294 491481
rect 157243 491409 157249 491469
rect 157283 491409 157294 491469
rect 157243 491397 157294 491409
rect 157384 491405 157418 491657
rect 156798 491233 156828 491397
rect 156865 491359 156957 491365
rect 156865 491325 156877 491359
rect 156945 491325 156957 491359
rect 156865 491319 156957 491325
rect 157141 491359 157233 491365
rect 157141 491325 157153 491359
rect 157221 491325 157233 491359
rect 157141 491319 157233 491325
rect 157264 491233 157294 491397
rect 143127 491191 157296 491233
rect 157254 491189 157296 491191
rect 147306 491085 147446 491097
rect 147306 491029 147346 491085
rect 147424 491029 147446 491085
rect 147306 490415 147446 491029
rect 158318 490600 159188 491657
rect 230433 490873 231381 491842
rect 327846 491762 327986 491774
rect 323888 491686 323972 491718
rect 323888 491644 323904 491686
rect 323958 491644 323972 491686
rect 323888 491556 323972 491644
rect 323888 491500 323896 491556
rect 323964 491500 323972 491556
rect 323888 491492 323972 491500
rect 327846 491706 327886 491762
rect 327964 491706 327986 491762
rect 247608 491127 249092 491157
rect 232818 491061 249092 491127
rect 327846 491092 327986 491706
rect 338790 491610 339590 492334
rect 418478 492100 418924 492104
rect 418118 492060 418924 492100
rect 418118 491900 418178 492060
rect 418338 491900 418924 492060
rect 419380 492016 419564 493280
rect 509380 492678 509564 493280
rect 509368 492592 510088 492678
rect 510002 492392 510088 492592
rect 510002 492328 510008 492392
rect 510080 492328 510088 492392
rect 510002 492302 510088 492328
rect 420030 492060 420570 492100
rect 419380 491924 419573 492016
rect 418118 491860 418924 491900
rect 418478 491854 418924 491860
rect 418723 491816 418923 491854
rect 419395 491844 419573 491924
rect 338790 491364 338860 491610
rect 339000 491364 339590 491610
rect 418821 491610 418851 491816
rect 419395 491784 419441 491844
rect 419535 491784 419573 491844
rect 420030 491900 420378 492060
rect 420538 491900 420570 492060
rect 509006 491996 512804 492050
rect 420030 491842 420570 491900
rect 508891 491843 508983 491849
rect 420073 491816 420273 491842
rect 419395 491750 419573 491784
rect 418821 491582 419971 491610
rect 418821 491443 418851 491582
rect 418890 491515 418982 491521
rect 418890 491481 418902 491515
rect 418970 491481 418982 491515
rect 418890 491475 418982 491481
rect 419166 491515 419258 491521
rect 419166 491481 419178 491515
rect 419246 491481 419258 491515
rect 419166 491475 419258 491481
rect 419015 491443 419049 491446
rect 418821 491431 418880 491443
rect 418821 491371 418840 491431
rect 418874 491371 418880 491431
rect 418821 491368 418880 491371
rect 338790 491278 339590 491364
rect 418834 491359 418880 491368
rect 418992 491431 419049 491443
rect 418992 491371 418998 491431
rect 419032 491412 419049 491431
rect 419101 491443 419137 491448
rect 419293 491443 419327 491582
rect 419101 491431 419156 491443
rect 419032 491371 419051 491412
rect 418992 491359 419051 491371
rect 418890 491321 418982 491327
rect 418890 491287 418902 491321
rect 418970 491287 418982 491321
rect 418890 491281 418982 491287
rect 418901 491244 418969 491281
rect 418901 491210 418923 491244
rect 418961 491210 418969 491244
rect 232698 490957 232790 490963
rect 232698 490923 232710 490957
rect 232778 490923 232790 490957
rect 232698 490917 232790 490923
rect 232823 490885 232863 491061
rect 232642 490873 232688 490885
rect 230433 490815 232648 490873
rect 230433 490798 231381 490815
rect 141258 488634 142348 488640
rect 143138 490215 147492 490415
rect 60798 488060 61758 488220
rect 143138 485815 143338 490215
rect 232484 490637 232526 490815
rect 232642 490813 232648 490815
rect 232682 490813 232688 490873
rect 232642 490801 232688 490813
rect 232800 490873 232863 490885
rect 232800 490813 232806 490873
rect 232840 490813 232863 490873
rect 232800 490801 232863 490813
rect 232823 490795 232863 490801
rect 232905 490885 232945 491061
rect 232974 490957 233066 490963
rect 232974 490923 232986 490957
rect 233054 490923 233066 490957
rect 232974 490917 233066 490923
rect 233250 490957 233342 490963
rect 233250 490923 233262 490957
rect 233330 490923 233342 490957
rect 233250 490917 233342 490923
rect 233099 490885 233129 490893
rect 232905 490873 232964 490885
rect 232905 490813 232924 490873
rect 232958 490813 232964 490873
rect 232905 490801 232964 490813
rect 233076 490873 233129 490885
rect 233076 490813 233082 490873
rect 233116 490813 233129 490873
rect 233076 490801 233129 490813
rect 232905 490797 232945 490801
rect 232698 490763 232790 490769
rect 232698 490729 232710 490763
rect 232778 490729 232790 490763
rect 232698 490723 232790 490729
rect 232974 490763 233066 490769
rect 232974 490729 232986 490763
rect 233054 490729 233066 490763
rect 232974 490723 233066 490729
rect 233099 490637 233129 490801
rect 233185 490885 233215 490893
rect 233381 490885 233421 491061
rect 233185 490873 233240 490885
rect 233185 490813 233200 490873
rect 233234 490813 233240 490873
rect 233185 490801 233240 490813
rect 233352 490873 233421 490885
rect 233352 490813 233358 490873
rect 233392 490813 233421 490873
rect 233352 490801 233421 490813
rect 233185 490637 233215 490801
rect 233381 490797 233421 490801
rect 233449 490885 233489 491061
rect 233526 490957 233618 490963
rect 233526 490923 233538 490957
rect 233606 490923 233618 490957
rect 233526 490917 233618 490923
rect 233802 490957 233894 490963
rect 233802 490923 233814 490957
rect 233882 490923 233894 490957
rect 233802 490917 233894 490923
rect 233653 490885 233683 490893
rect 233449 490873 233516 490885
rect 233449 490813 233476 490873
rect 233510 490813 233516 490873
rect 233449 490801 233516 490813
rect 233628 490873 233683 490885
rect 233628 490813 233634 490873
rect 233668 490813 233683 490873
rect 233628 490801 233683 490813
rect 233449 490797 233489 490801
rect 233250 490763 233342 490769
rect 233250 490729 233262 490763
rect 233330 490729 233342 490763
rect 233250 490723 233342 490729
rect 233526 490763 233618 490769
rect 233526 490729 233538 490763
rect 233606 490729 233618 490763
rect 233526 490723 233618 490729
rect 233653 490637 233683 490801
rect 233739 490885 233769 490893
rect 233929 490885 233969 491061
rect 233739 490873 233792 490885
rect 233739 490813 233752 490873
rect 233786 490813 233792 490873
rect 233739 490801 233792 490813
rect 233904 490873 233969 490885
rect 233904 490813 233910 490873
rect 233944 490813 233969 490873
rect 233904 490801 233969 490813
rect 233739 490637 233769 490801
rect 233929 490793 233969 490801
rect 234001 490885 234041 491061
rect 234078 490957 234170 490963
rect 234078 490923 234090 490957
rect 234158 490923 234170 490957
rect 234078 490917 234170 490923
rect 234354 490957 234446 490963
rect 234354 490923 234366 490957
rect 234434 490923 234446 490957
rect 234354 490917 234446 490923
rect 234201 490885 234231 490893
rect 234001 490873 234068 490885
rect 234001 490813 234028 490873
rect 234062 490813 234068 490873
rect 234001 490801 234068 490813
rect 234180 490873 234231 490885
rect 234180 490813 234186 490873
rect 234220 490813 234231 490873
rect 234180 490801 234231 490813
rect 234001 490797 234041 490801
rect 233802 490763 233894 490769
rect 233802 490729 233814 490763
rect 233882 490729 233894 490763
rect 233802 490723 233894 490729
rect 234078 490763 234170 490769
rect 234078 490729 234090 490763
rect 234158 490729 234170 490763
rect 234078 490723 234170 490729
rect 234201 490637 234231 490801
rect 234293 490885 234323 490891
rect 234481 490885 234521 491061
rect 234293 490873 234344 490885
rect 234293 490813 234304 490873
rect 234338 490813 234344 490873
rect 234293 490801 234344 490813
rect 234456 490873 234521 490885
rect 234456 490813 234462 490873
rect 234496 490813 234521 490873
rect 234456 490801 234521 490813
rect 234561 490885 234601 491061
rect 234630 490957 234722 490963
rect 234630 490923 234642 490957
rect 234710 490923 234722 490957
rect 234630 490917 234722 490923
rect 234906 490957 234998 490963
rect 234906 490923 234918 490957
rect 234986 490923 234998 490957
rect 234906 490917 234998 490923
rect 234751 490885 234781 490891
rect 234561 490873 234620 490885
rect 234561 490813 234580 490873
rect 234614 490813 234620 490873
rect 234561 490801 234620 490813
rect 234732 490873 234781 490885
rect 234732 490813 234738 490873
rect 234772 490813 234781 490873
rect 234732 490801 234781 490813
rect 234293 490637 234323 490801
rect 234354 490763 234446 490769
rect 234354 490729 234366 490763
rect 234434 490729 234446 490763
rect 234354 490723 234446 490729
rect 234630 490763 234722 490769
rect 234630 490729 234642 490763
rect 234710 490729 234722 490763
rect 234630 490723 234722 490729
rect 234751 490637 234781 490801
rect 234843 490885 234873 490889
rect 235035 490885 235075 491061
rect 234843 490873 234896 490885
rect 234843 490813 234856 490873
rect 234890 490813 234896 490873
rect 234843 490801 234896 490813
rect 235008 490873 235075 490885
rect 235008 490813 235014 490873
rect 235048 490813 235075 490873
rect 235008 490801 235075 490813
rect 234843 490637 234873 490801
rect 235035 490797 235075 490801
rect 235109 490885 235149 491061
rect 235182 490957 235274 490963
rect 235182 490923 235194 490957
rect 235262 490923 235274 490957
rect 235182 490917 235274 490923
rect 235458 490957 235550 490963
rect 235458 490923 235470 490957
rect 235538 490923 235550 490957
rect 235458 490917 235550 490923
rect 235307 490885 235337 490889
rect 235109 490873 235172 490885
rect 235109 490813 235132 490873
rect 235166 490813 235172 490873
rect 235109 490801 235172 490813
rect 235284 490873 235337 490885
rect 235284 490813 235290 490873
rect 235324 490813 235337 490873
rect 235284 490801 235337 490813
rect 235109 490799 235149 490801
rect 234906 490763 234998 490769
rect 234906 490729 234918 490763
rect 234986 490729 234998 490763
rect 234906 490723 234998 490729
rect 235182 490763 235274 490769
rect 235182 490729 235194 490763
rect 235262 490729 235274 490763
rect 235182 490723 235274 490729
rect 235307 490637 235337 490801
rect 235395 490885 235425 490887
rect 235587 490885 235627 491061
rect 235395 490873 235448 490885
rect 235395 490813 235408 490873
rect 235442 490813 235448 490873
rect 235395 490801 235448 490813
rect 235560 490873 235627 490885
rect 235560 490813 235566 490873
rect 235600 490813 235627 490873
rect 235560 490801 235627 490813
rect 235395 490637 235425 490801
rect 235587 490795 235627 490801
rect 235657 490885 235697 491061
rect 235734 490957 235826 490963
rect 235734 490923 235746 490957
rect 235814 490923 235826 490957
rect 235734 490917 235826 490923
rect 236010 490957 236102 490963
rect 236010 490923 236022 490957
rect 236090 490923 236102 490957
rect 236010 490917 236102 490923
rect 235857 490885 235887 490887
rect 235657 490873 235724 490885
rect 235657 490813 235684 490873
rect 235718 490813 235724 490873
rect 235657 490801 235724 490813
rect 235836 490873 235887 490885
rect 235836 490813 235842 490873
rect 235876 490813 235887 490873
rect 235836 490801 235887 490813
rect 235657 490799 235697 490801
rect 235458 490763 235550 490769
rect 235734 490767 235826 490769
rect 235458 490729 235470 490763
rect 235538 490729 235550 490763
rect 235731 490763 235826 490767
rect 235731 490734 235746 490763
rect 235458 490723 235550 490729
rect 235734 490729 235746 490734
rect 235814 490729 235826 490763
rect 235734 490723 235826 490729
rect 235857 490637 235887 490801
rect 235945 490885 235975 490887
rect 236135 490885 236175 491061
rect 235945 490873 236000 490885
rect 235945 490813 235960 490873
rect 235994 490813 236000 490873
rect 235945 490801 236000 490813
rect 236112 490873 236175 490885
rect 236112 490813 236118 490873
rect 236152 490813 236175 490873
rect 236112 490801 236175 490813
rect 235945 490637 235975 490801
rect 236135 490795 236175 490801
rect 236213 490885 236253 491061
rect 236286 490957 236378 490963
rect 236286 490923 236298 490957
rect 236366 490923 236378 490957
rect 236286 490917 236378 490923
rect 236562 490957 236654 490963
rect 236562 490923 236574 490957
rect 236642 490923 236654 490957
rect 236562 490917 236654 490923
rect 236409 490885 236439 490889
rect 236213 490873 236276 490885
rect 236213 490813 236236 490873
rect 236270 490813 236276 490873
rect 236213 490801 236276 490813
rect 236388 490873 236439 490885
rect 236388 490813 236394 490873
rect 236428 490813 236439 490873
rect 236388 490801 236439 490813
rect 236213 490799 236253 490801
rect 236010 490763 236102 490769
rect 236010 490729 236022 490763
rect 236090 490729 236102 490763
rect 236010 490723 236102 490729
rect 236286 490763 236378 490769
rect 236286 490729 236298 490763
rect 236366 490729 236378 490763
rect 236286 490723 236378 490729
rect 236409 490637 236439 490801
rect 236497 490885 236527 490889
rect 236689 490885 236729 491061
rect 236497 490873 236552 490885
rect 236497 490813 236512 490873
rect 236546 490813 236552 490873
rect 236497 490801 236552 490813
rect 236664 490873 236729 490885
rect 236664 490813 236670 490873
rect 236704 490813 236729 490873
rect 236664 490801 236729 490813
rect 236497 490637 236527 490801
rect 236689 490787 236729 490801
rect 236767 490885 236807 491061
rect 236838 490957 236930 490963
rect 236838 490923 236850 490957
rect 236918 490923 236930 490957
rect 236838 490917 236930 490923
rect 237114 490957 237206 490963
rect 237114 490923 237126 490957
rect 237194 490923 237206 490957
rect 237114 490917 237206 490923
rect 236961 490885 236991 490889
rect 236767 490873 236828 490885
rect 236767 490813 236788 490873
rect 236822 490813 236828 490873
rect 236767 490801 236828 490813
rect 236940 490873 236991 490885
rect 236940 490813 236946 490873
rect 236980 490813 236991 490873
rect 236940 490801 236991 490813
rect 236767 490795 236807 490801
rect 236562 490763 236654 490769
rect 236562 490729 236574 490763
rect 236642 490729 236654 490763
rect 236562 490723 236654 490729
rect 236838 490763 236930 490769
rect 236838 490729 236850 490763
rect 236918 490729 236930 490763
rect 236838 490723 236930 490729
rect 236961 490637 236991 490801
rect 237053 490885 237083 490889
rect 237245 490885 237285 491061
rect 237053 490873 237104 490885
rect 237053 490813 237064 490873
rect 237098 490813 237104 490873
rect 237053 490801 237104 490813
rect 237216 490873 237285 490885
rect 237216 490813 237222 490873
rect 237256 490813 237285 490873
rect 237216 490801 237285 490813
rect 237319 490885 237359 491061
rect 237390 490957 237482 490963
rect 237390 490923 237402 490957
rect 237470 490923 237482 490957
rect 237390 490917 237482 490923
rect 237666 490957 237758 490963
rect 237666 490923 237678 490957
rect 237746 490923 237758 490957
rect 237666 490917 237758 490923
rect 237515 490885 237545 490899
rect 237319 490873 237380 490885
rect 237319 490813 237340 490873
rect 237374 490813 237380 490873
rect 237319 490801 237380 490813
rect 237492 490873 237545 490885
rect 237492 490813 237498 490873
rect 237532 490813 237545 490873
rect 237492 490801 237545 490813
rect 237053 490637 237083 490801
rect 237245 490797 237285 490801
rect 237114 490763 237206 490769
rect 237114 490729 237126 490763
rect 237194 490729 237206 490763
rect 237114 490723 237206 490729
rect 237390 490763 237482 490769
rect 237390 490729 237402 490763
rect 237470 490729 237482 490763
rect 237390 490723 237482 490729
rect 237515 490637 237545 490801
rect 237601 490885 237631 490897
rect 237789 490885 237823 491061
rect 237601 490873 237656 490885
rect 237601 490813 237616 490873
rect 237650 490813 237656 490873
rect 237601 490801 237656 490813
rect 237768 490873 237823 490885
rect 237768 490813 237774 490873
rect 237808 490813 237823 490873
rect 237768 490801 237823 490813
rect 237601 490637 237631 490801
rect 237789 490797 237823 490801
rect 237879 490885 237913 491061
rect 237942 490957 238034 490963
rect 237942 490923 237954 490957
rect 238022 490923 238034 490957
rect 237942 490917 238034 490923
rect 238218 490957 238310 490963
rect 238218 490923 238230 490957
rect 238298 490923 238310 490957
rect 238218 490917 238310 490923
rect 238069 490885 238099 490895
rect 237879 490873 237932 490885
rect 237879 490813 237892 490873
rect 237926 490813 237932 490873
rect 237879 490801 237932 490813
rect 238044 490873 238099 490885
rect 238044 490813 238050 490873
rect 238084 490813 238099 490873
rect 238044 490801 238099 490813
rect 237879 490797 237913 490801
rect 237666 490763 237758 490769
rect 237666 490729 237678 490763
rect 237746 490729 237758 490763
rect 237666 490723 237758 490729
rect 237942 490763 238034 490769
rect 237942 490729 237954 490763
rect 238022 490729 238034 490763
rect 237942 490723 238034 490729
rect 238069 490637 238099 490801
rect 238155 490885 238185 490895
rect 238345 490885 238379 491061
rect 238155 490873 238208 490885
rect 238155 490813 238168 490873
rect 238202 490813 238208 490873
rect 238155 490801 238208 490813
rect 238320 490873 238379 490885
rect 238320 490813 238326 490873
rect 238360 490813 238379 490873
rect 238320 490801 238379 490813
rect 238429 490885 238463 491061
rect 238494 490957 238586 490963
rect 238494 490923 238506 490957
rect 238574 490923 238586 490957
rect 238494 490917 238586 490923
rect 238621 490885 238655 490899
rect 238429 490873 238484 490885
rect 238429 490813 238444 490873
rect 238478 490813 238484 490873
rect 238429 490801 238484 490813
rect 238596 490873 238655 490885
rect 238596 490813 238602 490873
rect 238636 490813 238655 490873
rect 238596 490801 238655 490813
rect 238155 490637 238185 490801
rect 238345 490797 238379 490801
rect 238218 490763 238310 490769
rect 238218 490729 238230 490763
rect 238298 490729 238310 490763
rect 238218 490723 238310 490729
rect 238494 490763 238586 490769
rect 238494 490729 238506 490763
rect 238574 490729 238586 490763
rect 238494 490723 238586 490729
rect 238621 490637 238655 490801
rect 238703 490885 238737 491061
rect 238770 490957 238862 490963
rect 238770 490923 238782 490957
rect 238850 490923 238862 490957
rect 238770 490917 238862 490923
rect 239046 490957 239138 490963
rect 239046 490923 239058 490957
rect 239126 490923 239138 490957
rect 239046 490917 239138 490923
rect 238895 490885 238925 490897
rect 238703 490873 238760 490885
rect 238703 490813 238720 490873
rect 238754 490813 238760 490873
rect 238703 490801 238760 490813
rect 238872 490873 238925 490885
rect 238872 490813 238878 490873
rect 238912 490813 238925 490873
rect 238872 490801 238925 490813
rect 238703 490799 238737 490801
rect 238770 490763 238862 490769
rect 238770 490729 238782 490763
rect 238850 490729 238862 490763
rect 238770 490723 238862 490729
rect 238895 490637 238925 490801
rect 238983 490885 239013 490899
rect 239173 490885 239207 491061
rect 238983 490873 239036 490885
rect 238983 490813 238996 490873
rect 239030 490813 239036 490873
rect 238983 490801 239036 490813
rect 239148 490873 239207 490885
rect 239148 490813 239154 490873
rect 239188 490813 239207 490873
rect 239148 490801 239207 490813
rect 239259 490885 239293 491061
rect 239331 490999 239546 491009
rect 239331 490963 239461 490999
rect 239322 490957 239461 490963
rect 239322 490923 239334 490957
rect 239402 490939 239461 490957
rect 239521 490939 239546 490999
rect 239402 490929 239546 490939
rect 239598 490957 239690 490963
rect 239402 490923 239414 490929
rect 239322 490917 239414 490923
rect 239598 490923 239610 490957
rect 239678 490923 239690 490957
rect 239598 490917 239690 490923
rect 239443 490885 239473 490899
rect 239259 490873 239312 490885
rect 239259 490813 239272 490873
rect 239306 490813 239312 490873
rect 239259 490801 239312 490813
rect 239424 490873 239473 490885
rect 239424 490813 239430 490873
rect 239464 490813 239473 490873
rect 239424 490801 239473 490813
rect 238983 490637 239013 490801
rect 239259 490795 239293 490801
rect 239046 490763 239138 490769
rect 239046 490729 239058 490763
rect 239126 490729 239138 490763
rect 239322 490763 239414 490769
rect 239322 490744 239334 490763
rect 239046 490723 239138 490729
rect 239186 490739 239334 490744
rect 239186 490684 239196 490739
rect 239261 490729 239334 490739
rect 239402 490729 239414 490763
rect 239261 490723 239414 490729
rect 239261 490694 239401 490723
rect 239261 490684 239271 490694
rect 239186 490679 239271 490684
rect 239443 490637 239473 490801
rect 239535 490885 239565 490899
rect 239725 490885 239759 491061
rect 239535 490873 239588 490885
rect 239535 490813 239548 490873
rect 239582 490813 239588 490873
rect 239535 490801 239588 490813
rect 239700 490873 239759 490885
rect 239700 490813 239706 490873
rect 239740 490813 239759 490873
rect 239700 490803 239759 490813
rect 239811 490885 239845 491061
rect 239874 490957 239966 490963
rect 239874 490923 239886 490957
rect 239954 490923 239966 490957
rect 239874 490917 239966 490923
rect 240150 490957 240242 490963
rect 240150 490923 240162 490957
rect 240230 490923 240242 490957
rect 240150 490917 240242 490923
rect 239997 490885 240027 490899
rect 239811 490873 239864 490885
rect 239811 490813 239824 490873
rect 239858 490813 239864 490873
rect 239700 490801 239746 490803
rect 239811 490801 239864 490813
rect 239976 490873 240027 490885
rect 239976 490813 239982 490873
rect 240016 490813 240027 490873
rect 239976 490801 240027 490813
rect 239535 490637 239565 490801
rect 239811 490799 239845 490801
rect 239598 490763 239690 490769
rect 239598 490729 239610 490763
rect 239678 490729 239690 490763
rect 239598 490723 239690 490729
rect 239874 490763 239966 490769
rect 239874 490729 239886 490763
rect 239954 490729 239966 490763
rect 239874 490723 239966 490729
rect 239997 490637 240027 490801
rect 240089 490885 240119 490899
rect 240275 490885 240309 491061
rect 240089 490873 240140 490885
rect 240089 490813 240100 490873
rect 240134 490813 240140 490873
rect 240089 490801 240140 490813
rect 240252 490873 240309 490885
rect 240252 490813 240258 490873
rect 240292 490813 240309 490873
rect 240252 490801 240309 490813
rect 240089 490637 240119 490801
rect 240275 490799 240309 490801
rect 240363 490885 240397 491061
rect 240426 490957 240518 490963
rect 240426 490923 240438 490957
rect 240506 490923 240518 490957
rect 240426 490917 240518 490923
rect 240702 490957 240794 490963
rect 240702 490923 240714 490957
rect 240782 490923 240794 490957
rect 240702 490917 240794 490923
rect 240549 490885 240579 490899
rect 240363 490873 240416 490885
rect 240363 490813 240376 490873
rect 240410 490813 240416 490873
rect 240363 490801 240416 490813
rect 240528 490873 240579 490885
rect 240528 490813 240534 490873
rect 240568 490813 240579 490873
rect 240528 490801 240579 490813
rect 240363 490797 240397 490801
rect 240150 490763 240242 490769
rect 240150 490729 240162 490763
rect 240230 490729 240242 490763
rect 240150 490723 240242 490729
rect 240426 490763 240518 490769
rect 240426 490729 240438 490763
rect 240506 490729 240518 490763
rect 240426 490723 240518 490729
rect 240549 490637 240579 490801
rect 240635 490885 240665 490899
rect 240831 490885 240865 491061
rect 240635 490873 240692 490885
rect 240635 490813 240652 490873
rect 240686 490813 240692 490873
rect 240635 490801 240692 490813
rect 240804 490873 240865 490885
rect 240804 490813 240810 490873
rect 240844 490813 240865 490873
rect 240804 490801 240865 490813
rect 240635 490637 240665 490801
rect 240831 490793 240865 490801
rect 240913 490885 240947 491061
rect 240978 490957 241070 490963
rect 240978 490923 240990 490957
rect 241058 490923 241070 490957
rect 240978 490917 241070 490923
rect 241254 490957 241346 490963
rect 241254 490923 241266 490957
rect 241334 490923 241346 490957
rect 241254 490917 241346 490923
rect 241103 490885 241133 490899
rect 240913 490873 240968 490885
rect 240913 490813 240928 490873
rect 240962 490813 240968 490873
rect 240913 490801 240968 490813
rect 241080 490873 241133 490885
rect 241080 490813 241086 490873
rect 241120 490813 241133 490873
rect 241080 490801 241133 490813
rect 240913 490799 240947 490801
rect 240702 490763 240794 490769
rect 240702 490729 240714 490763
rect 240782 490729 240794 490763
rect 240702 490723 240794 490729
rect 240978 490763 241070 490769
rect 240978 490729 240990 490763
rect 241058 490729 241070 490763
rect 240978 490723 241070 490729
rect 241103 490637 241133 490801
rect 241191 490885 241221 490897
rect 241385 490885 241419 491061
rect 241191 490873 241244 490885
rect 241191 490813 241204 490873
rect 241238 490813 241244 490873
rect 241191 490801 241244 490813
rect 241356 490873 241419 490885
rect 241356 490813 241362 490873
rect 241396 490813 241419 490873
rect 241356 490801 241419 490813
rect 241191 490637 241221 490801
rect 241385 490797 241419 490801
rect 241463 490885 241497 491061
rect 241530 490957 241622 490963
rect 241530 490923 241542 490957
rect 241610 490923 241622 490957
rect 241530 490917 241622 490923
rect 241806 490957 241898 490963
rect 241806 490923 241818 490957
rect 241886 490923 241898 490957
rect 241806 490917 241898 490923
rect 241655 490885 241685 490901
rect 241463 490873 241520 490885
rect 241463 490813 241480 490873
rect 241514 490813 241520 490873
rect 241463 490801 241520 490813
rect 241632 490873 241685 490885
rect 241632 490813 241638 490873
rect 241672 490813 241685 490873
rect 241632 490801 241685 490813
rect 241463 490799 241497 490801
rect 241254 490763 241346 490769
rect 241254 490729 241266 490763
rect 241334 490729 241346 490763
rect 241254 490723 241346 490729
rect 241530 490763 241622 490769
rect 241530 490729 241542 490763
rect 241610 490729 241622 490763
rect 241530 490723 241622 490729
rect 241655 490637 241685 490801
rect 241743 490885 241773 490901
rect 241941 490885 241975 491061
rect 241743 490873 241796 490885
rect 241743 490813 241756 490873
rect 241790 490813 241796 490873
rect 241743 490801 241796 490813
rect 241908 490873 241975 490885
rect 241908 490813 241914 490873
rect 241948 490813 241975 490873
rect 241908 490801 241975 490813
rect 241743 490637 241773 490801
rect 241941 490789 241975 490801
rect 242015 490885 242049 491061
rect 242082 490957 242174 490963
rect 242082 490923 242094 490957
rect 242162 490923 242174 490957
rect 242082 490917 242174 490923
rect 242358 490957 242450 490963
rect 242358 490923 242370 490957
rect 242438 490923 242450 490957
rect 242358 490917 242450 490923
rect 242205 490885 242235 490903
rect 242015 490873 242072 490885
rect 242015 490813 242032 490873
rect 242066 490813 242072 490873
rect 242015 490801 242072 490813
rect 242184 490873 242235 490885
rect 242184 490813 242190 490873
rect 242224 490813 242235 490873
rect 242184 490801 242235 490813
rect 242015 490793 242049 490801
rect 241806 490763 241898 490769
rect 241806 490729 241818 490763
rect 241886 490729 241898 490763
rect 241806 490723 241898 490729
rect 242082 490763 242174 490769
rect 242082 490729 242094 490763
rect 242162 490729 242174 490763
rect 242082 490723 242174 490729
rect 242205 490637 242235 490801
rect 242293 490885 242323 490901
rect 242485 490885 242519 491061
rect 242293 490873 242348 490885
rect 242293 490813 242308 490873
rect 242342 490813 242348 490873
rect 242293 490801 242348 490813
rect 242460 490873 242519 490885
rect 242460 490813 242466 490873
rect 242500 490813 242519 490873
rect 242460 490801 242519 490813
rect 242293 490637 242323 490801
rect 242485 490789 242519 490801
rect 242565 490885 242599 491061
rect 242634 490957 242726 490963
rect 242634 490923 242646 490957
rect 242714 490923 242726 490957
rect 242634 490917 242726 490923
rect 242910 490957 243002 490963
rect 242910 490923 242922 490957
rect 242990 490923 243002 490957
rect 242910 490917 243002 490923
rect 242757 490885 242787 490901
rect 242565 490873 242624 490885
rect 242565 490813 242584 490873
rect 242618 490813 242624 490873
rect 242565 490801 242624 490813
rect 242736 490873 242787 490885
rect 242736 490813 242742 490873
rect 242776 490813 242787 490873
rect 242736 490801 242787 490813
rect 242565 490787 242599 490801
rect 242358 490763 242450 490769
rect 242358 490729 242370 490763
rect 242438 490729 242450 490763
rect 242358 490723 242450 490729
rect 242634 490763 242726 490769
rect 242634 490729 242646 490763
rect 242714 490729 242726 490763
rect 242634 490723 242726 490729
rect 242757 490637 242787 490801
rect 242845 490885 242875 490903
rect 243041 490885 243075 491061
rect 242845 490873 242900 490885
rect 242845 490813 242860 490873
rect 242894 490813 242900 490873
rect 242845 490801 242900 490813
rect 243012 490873 243075 490885
rect 243012 490813 243018 490873
rect 243052 490813 243075 490873
rect 243012 490801 243075 490813
rect 242845 490637 242875 490801
rect 243041 490789 243075 490801
rect 243115 490885 243149 491061
rect 243186 490957 243278 490963
rect 243186 490923 243198 490957
rect 243266 490923 243278 490957
rect 243186 490917 243278 490923
rect 243462 490957 243554 490963
rect 243462 490923 243474 490957
rect 243542 490923 243554 490957
rect 243462 490917 243554 490923
rect 243309 490885 243339 490901
rect 243115 490873 243176 490885
rect 243115 490813 243136 490873
rect 243170 490813 243176 490873
rect 243115 490801 243176 490813
rect 243288 490873 243339 490885
rect 243288 490813 243294 490873
rect 243328 490813 243339 490873
rect 243288 490801 243339 490813
rect 243115 490787 243149 490801
rect 242910 490763 243002 490769
rect 242910 490729 242922 490763
rect 242990 490729 243002 490763
rect 242910 490723 243002 490729
rect 243186 490763 243278 490769
rect 243186 490729 243198 490763
rect 243266 490729 243278 490763
rect 243186 490723 243278 490729
rect 243309 490637 243339 490801
rect 243399 490885 243429 490903
rect 243591 490885 243625 491061
rect 243399 490873 243452 490885
rect 243399 490813 243412 490873
rect 243446 490813 243452 490873
rect 243399 490801 243452 490813
rect 243564 490873 243625 490885
rect 243564 490813 243570 490873
rect 243604 490813 243625 490873
rect 243564 490801 243625 490813
rect 243399 490637 243429 490801
rect 243591 490791 243625 490801
rect 243667 490885 243701 491061
rect 243738 490957 243830 490963
rect 243738 490923 243750 490957
rect 243818 490923 243830 490957
rect 243738 490917 243830 490923
rect 244014 490957 244106 490963
rect 244014 490923 244026 490957
rect 244094 490923 244106 490957
rect 244014 490917 244106 490923
rect 243861 490885 243891 490901
rect 243667 490873 243728 490885
rect 243667 490813 243688 490873
rect 243722 490813 243728 490873
rect 243667 490801 243728 490813
rect 243840 490873 243891 490885
rect 243840 490813 243846 490873
rect 243880 490813 243891 490873
rect 243840 490801 243891 490813
rect 243667 490791 243701 490801
rect 243462 490763 243554 490769
rect 243462 490729 243474 490763
rect 243542 490729 243554 490763
rect 243462 490723 243554 490729
rect 243738 490763 243830 490769
rect 243738 490729 243750 490763
rect 243818 490729 243830 490763
rect 243738 490723 243830 490729
rect 243861 490637 243891 490801
rect 243951 490885 243981 490903
rect 244141 490885 244175 491061
rect 243951 490873 244004 490885
rect 243951 490813 243964 490873
rect 243998 490813 244004 490873
rect 243951 490801 244004 490813
rect 244116 490873 244175 490885
rect 244116 490813 244122 490873
rect 244156 490813 244175 490873
rect 244116 490801 244175 490813
rect 243951 490637 243981 490801
rect 244141 490795 244175 490801
rect 244223 490885 244257 491061
rect 244290 490957 244382 490963
rect 244290 490923 244302 490957
rect 244370 490923 244382 490957
rect 244290 490917 244382 490923
rect 244566 490957 244658 490963
rect 244566 490923 244578 490957
rect 244646 490923 244658 490957
rect 244566 490917 244658 490923
rect 244415 490885 244445 490907
rect 244223 490873 244280 490885
rect 244223 490813 244240 490873
rect 244274 490813 244280 490873
rect 244223 490801 244280 490813
rect 244392 490873 244445 490885
rect 244392 490813 244398 490873
rect 244432 490813 244445 490873
rect 244392 490801 244445 490813
rect 244223 490793 244257 490801
rect 244014 490763 244106 490769
rect 244014 490729 244026 490763
rect 244094 490729 244106 490763
rect 244014 490723 244106 490729
rect 244290 490763 244382 490769
rect 244290 490729 244302 490763
rect 244370 490729 244382 490763
rect 244290 490723 244382 490729
rect 244415 490637 244445 490801
rect 244505 490885 244535 490909
rect 244693 490885 244727 491061
rect 244505 490873 244556 490885
rect 244505 490813 244516 490873
rect 244550 490813 244556 490873
rect 244505 490801 244556 490813
rect 244668 490873 244727 490885
rect 244668 490813 244674 490873
rect 244708 490813 244727 490873
rect 244668 490801 244727 490813
rect 244771 490885 244805 491061
rect 244842 490957 244934 490963
rect 244842 490923 244854 490957
rect 244922 490923 244934 490957
rect 244842 490917 244934 490923
rect 245118 490957 245210 490963
rect 245118 490923 245130 490957
rect 245198 490923 245210 490957
rect 245118 490917 245210 490923
rect 244969 490885 244999 490909
rect 244771 490873 244832 490885
rect 244771 490813 244792 490873
rect 244826 490813 244832 490873
rect 244771 490801 244832 490813
rect 244944 490873 244999 490885
rect 244944 490813 244950 490873
rect 244984 490813 244999 490873
rect 244944 490801 244999 490813
rect 244505 490637 244535 490801
rect 244693 490799 244727 490801
rect 244566 490763 244658 490769
rect 244566 490729 244578 490763
rect 244646 490729 244658 490763
rect 244566 490723 244658 490729
rect 244842 490763 244934 490769
rect 244842 490729 244854 490763
rect 244922 490729 244934 490763
rect 244842 490723 244934 490729
rect 244969 490637 244999 490801
rect 245055 490885 245085 490913
rect 245243 490885 245277 491061
rect 245055 490873 245108 490885
rect 245055 490813 245068 490873
rect 245102 490813 245108 490873
rect 245055 490801 245108 490813
rect 245220 490873 245277 490885
rect 245220 490813 245226 490873
rect 245260 490813 245277 490873
rect 245220 490801 245277 490813
rect 245055 490637 245085 490801
rect 245243 490797 245277 490801
rect 245327 490885 245361 491061
rect 245394 490957 245486 490963
rect 245394 490923 245406 490957
rect 245474 490923 245486 490957
rect 245394 490917 245486 490923
rect 245670 490957 245762 490963
rect 245670 490923 245682 490957
rect 245750 490923 245762 490957
rect 245670 490917 245762 490923
rect 245515 490885 245545 490899
rect 245327 490873 245384 490885
rect 245327 490813 245344 490873
rect 245378 490813 245384 490873
rect 245327 490801 245384 490813
rect 245496 490873 245545 490885
rect 245496 490813 245502 490873
rect 245536 490813 245545 490873
rect 245496 490801 245545 490813
rect 245327 490795 245361 490801
rect 245118 490763 245210 490769
rect 245118 490729 245130 490763
rect 245198 490729 245210 490763
rect 245118 490723 245210 490729
rect 245394 490763 245486 490769
rect 245394 490729 245406 490763
rect 245474 490729 245486 490763
rect 245394 490723 245486 490729
rect 245515 490637 245545 490801
rect 245607 490885 245637 490897
rect 245795 490885 245829 491061
rect 245607 490873 245660 490885
rect 245607 490813 245620 490873
rect 245654 490813 245660 490873
rect 245607 490801 245660 490813
rect 245772 490873 245829 490885
rect 245772 490813 245778 490873
rect 245812 490813 245829 490873
rect 245772 490801 245829 490813
rect 245607 490637 245637 490801
rect 245795 490797 245829 490801
rect 245879 490885 245913 491061
rect 245946 490957 246038 490963
rect 245946 490923 245958 490957
rect 246026 490923 246038 490957
rect 245946 490917 246038 490923
rect 246222 490957 246314 490963
rect 246222 490923 246234 490957
rect 246302 490923 246314 490957
rect 246222 490917 246314 490923
rect 246071 490885 246101 490899
rect 245879 490873 245936 490885
rect 245879 490813 245896 490873
rect 245930 490813 245936 490873
rect 245879 490801 245936 490813
rect 246048 490873 246101 490885
rect 246048 490813 246054 490873
rect 246088 490813 246101 490873
rect 246048 490801 246101 490813
rect 245879 490799 245913 490801
rect 245670 490763 245762 490769
rect 245670 490729 245682 490763
rect 245750 490729 245762 490763
rect 245670 490723 245762 490729
rect 245946 490763 246038 490769
rect 245946 490729 245958 490763
rect 246026 490729 246038 490763
rect 245946 490723 246038 490729
rect 246071 490637 246101 490801
rect 246155 490885 246185 490899
rect 246349 490885 246383 491061
rect 246155 490873 246212 490885
rect 246155 490813 246172 490873
rect 246206 490813 246212 490873
rect 246155 490801 246212 490813
rect 246324 490873 246383 490885
rect 246324 490813 246330 490873
rect 246364 490813 246383 490873
rect 246324 490803 246383 490813
rect 246427 490885 246461 491061
rect 246498 490957 246590 490963
rect 246498 490923 246510 490957
rect 246578 490923 246590 490957
rect 246498 490917 246590 490923
rect 246621 490885 246651 490899
rect 246427 490873 246488 490885
rect 246427 490813 246448 490873
rect 246482 490813 246488 490873
rect 246324 490801 246370 490803
rect 246427 490801 246488 490813
rect 246600 490873 246651 490885
rect 246600 490813 246606 490873
rect 246640 490813 246651 490873
rect 246600 490801 246651 490813
rect 246741 490809 246775 491061
rect 246155 490637 246185 490801
rect 246222 490763 246314 490769
rect 246222 490729 246234 490763
rect 246302 490729 246314 490763
rect 246222 490723 246314 490729
rect 246498 490763 246590 490769
rect 246498 490729 246510 490763
rect 246578 490729 246590 490763
rect 246498 490723 246590 490729
rect 246621 490637 246651 490801
rect 232484 490595 246653 490637
rect 246611 490593 246653 490595
rect 236663 490489 236803 490501
rect 236663 490433 236703 490489
rect 236781 490433 236803 490489
rect 236663 489819 236803 490433
rect 247591 490134 249092 491061
rect 158318 489724 159188 489730
rect 233035 489619 236849 489819
rect 233035 487388 233235 489619
rect 322870 490892 328032 491092
rect 418901 491066 418969 491210
rect 419015 491175 419051 491359
rect 419101 491371 419116 491431
rect 419150 491371 419156 491431
rect 419101 491359 419156 491371
rect 419268 491431 419327 491443
rect 419268 491371 419274 491431
rect 419308 491371 419327 491431
rect 419268 491359 419327 491371
rect 419101 491175 419137 491359
rect 419293 491340 419327 491359
rect 419371 491443 419405 491582
rect 419437 491542 419539 491550
rect 419437 491484 419445 491542
rect 419531 491484 419539 491542
rect 419437 491481 419454 491484
rect 419522 491481 419539 491484
rect 419437 491476 419539 491481
rect 419718 491515 419810 491521
rect 419718 491481 419730 491515
rect 419798 491481 419810 491515
rect 419442 491475 419534 491476
rect 419718 491475 419810 491481
rect 419573 491443 419611 491444
rect 419851 491443 419885 491582
rect 419371 491431 419432 491443
rect 419371 491371 419392 491431
rect 419426 491371 419432 491431
rect 419371 491359 419432 491371
rect 419544 491431 419611 491443
rect 419662 491442 419708 491443
rect 419544 491371 419550 491431
rect 419584 491371 419611 491431
rect 419544 491359 419611 491371
rect 419371 491338 419405 491359
rect 419166 491321 419258 491327
rect 419442 491326 419534 491327
rect 419166 491287 419178 491321
rect 419246 491287 419258 491321
rect 419166 491281 419258 491287
rect 419437 491321 419539 491326
rect 419437 491318 419454 491321
rect 419522 491318 419539 491321
rect 419437 491260 419445 491318
rect 419531 491260 419539 491318
rect 419437 491252 419539 491260
rect 419015 491174 419295 491175
rect 419573 491174 419611 491359
rect 419647 491431 419708 491442
rect 419647 491371 419668 491431
rect 419702 491371 419708 491431
rect 419647 491359 419708 491371
rect 419820 491431 419885 491443
rect 419820 491371 419826 491431
rect 419860 491371 419885 491431
rect 419820 491359 419885 491371
rect 419647 491174 419685 491359
rect 419851 491340 419885 491359
rect 419921 491443 419955 491582
rect 419994 491515 420086 491521
rect 419994 491481 420006 491515
rect 420074 491481 420086 491515
rect 419994 491475 420086 491481
rect 420237 491444 420271 491816
rect 507964 491786 508164 491834
rect 508891 491809 508903 491843
rect 508971 491809 508983 491843
rect 508891 491803 508983 491809
rect 507964 491684 507996 491786
rect 508146 491684 508164 491786
rect 507964 491634 508164 491684
rect 508828 491771 508860 491788
rect 509012 491771 509042 491996
rect 508828 491759 508881 491771
rect 508828 491699 508841 491759
rect 508875 491699 508881 491759
rect 508828 491687 508881 491699
rect 508993 491759 509042 491771
rect 508993 491699 508999 491759
rect 509033 491699 509042 491759
rect 508993 491687 509042 491699
rect 420117 491443 420271 491444
rect 419921 491431 419984 491443
rect 419921 491371 419944 491431
rect 419978 491371 419984 491431
rect 419921 491359 419984 491371
rect 420096 491434 420271 491443
rect 508039 491434 508085 491634
rect 508828 491434 508860 491687
rect 509012 491666 509042 491687
rect 509102 491771 509132 491996
rect 509167 491843 509259 491849
rect 509167 491809 509179 491843
rect 509247 491809 509259 491843
rect 509167 491803 509259 491809
rect 509443 491843 509535 491849
rect 509443 491809 509455 491843
rect 509523 491809 509535 491843
rect 509443 491803 509535 491809
rect 509294 491771 509326 491790
rect 509102 491759 509157 491771
rect 509102 491699 509117 491759
rect 509151 491699 509157 491759
rect 509102 491687 509157 491699
rect 509269 491759 509326 491771
rect 509269 491699 509275 491759
rect 509309 491699 509326 491759
rect 509269 491687 509326 491699
rect 509102 491666 509132 491687
rect 508891 491649 508983 491655
rect 508891 491615 508903 491649
rect 508971 491615 508983 491649
rect 508891 491609 508983 491615
rect 509167 491649 509259 491655
rect 509167 491615 509179 491649
rect 509247 491615 509259 491649
rect 509167 491609 509259 491615
rect 509294 491434 509326 491687
rect 509376 491771 509408 491790
rect 509564 491771 509594 491996
rect 509376 491759 509433 491771
rect 509376 491699 509393 491759
rect 509427 491699 509433 491759
rect 509376 491687 509433 491699
rect 509545 491759 509594 491771
rect 509545 491699 509551 491759
rect 509585 491699 509594 491759
rect 509545 491687 509594 491699
rect 509376 491434 509408 491687
rect 509564 491668 509594 491687
rect 509654 491771 509684 491996
rect 510006 491872 510086 491882
rect 510006 491849 510008 491872
rect 509719 491843 509811 491849
rect 509719 491809 509731 491843
rect 509799 491809 509811 491843
rect 509719 491803 509811 491809
rect 509995 491843 510008 491849
rect 510076 491849 510086 491872
rect 509995 491809 510007 491843
rect 510076 491816 510087 491849
rect 510075 491809 510087 491816
rect 509995 491803 510087 491809
rect 509846 491771 509878 491790
rect 509654 491759 509709 491771
rect 509654 491699 509669 491759
rect 509703 491699 509709 491759
rect 509654 491687 509709 491699
rect 509821 491759 509878 491771
rect 509821 491699 509827 491759
rect 509861 491699 509878 491759
rect 509821 491687 509878 491699
rect 509654 491666 509684 491687
rect 509443 491649 509535 491655
rect 509443 491615 509455 491649
rect 509523 491615 509535 491649
rect 509443 491609 509535 491615
rect 509719 491649 509811 491655
rect 509719 491615 509731 491649
rect 509799 491615 509811 491649
rect 509719 491609 509811 491615
rect 509846 491434 509878 491687
rect 509934 491771 509966 491788
rect 510118 491771 510148 491996
rect 509934 491759 509985 491771
rect 509934 491699 509945 491759
rect 509979 491699 509985 491759
rect 509934 491687 509985 491699
rect 510097 491759 510148 491771
rect 510097 491699 510103 491759
rect 510137 491699 510148 491759
rect 510097 491687 510148 491699
rect 509934 491434 509966 491687
rect 510118 491662 510148 491687
rect 510208 491771 510238 491996
rect 510271 491843 510363 491849
rect 510271 491809 510283 491843
rect 510351 491809 510363 491843
rect 510271 491803 510363 491809
rect 510547 491843 510639 491849
rect 510547 491809 510559 491843
rect 510627 491809 510639 491843
rect 510547 491803 510639 491809
rect 510394 491771 510426 491790
rect 510208 491759 510261 491771
rect 510208 491699 510221 491759
rect 510255 491699 510261 491759
rect 510208 491687 510261 491699
rect 510373 491759 510426 491771
rect 510373 491699 510379 491759
rect 510413 491699 510426 491759
rect 510373 491687 510426 491699
rect 510208 491660 510238 491687
rect 510000 491655 510080 491656
rect 509995 491649 510087 491655
rect 509995 491615 510007 491649
rect 510075 491642 510087 491649
rect 509995 491609 510008 491615
rect 510000 491586 510008 491609
rect 510076 491609 510087 491642
rect 510271 491649 510363 491655
rect 510271 491615 510283 491649
rect 510351 491615 510363 491649
rect 510271 491609 510363 491615
rect 510076 491586 510080 491609
rect 510000 491578 510080 491586
rect 510394 491434 510426 491687
rect 510482 491771 510514 491788
rect 510668 491771 510698 491996
rect 510482 491759 510537 491771
rect 510482 491699 510497 491759
rect 510531 491699 510537 491759
rect 510482 491687 510537 491699
rect 510649 491759 510698 491771
rect 510649 491699 510655 491759
rect 510689 491699 510698 491759
rect 510649 491687 510698 491699
rect 510482 491434 510514 491687
rect 510668 491672 510698 491687
rect 510758 491771 510788 491996
rect 510823 491843 510915 491849
rect 510823 491809 510835 491843
rect 510903 491809 510915 491843
rect 510823 491803 510915 491809
rect 511099 491843 511191 491849
rect 511099 491809 511111 491843
rect 511179 491809 511191 491843
rect 511099 491803 511191 491809
rect 510946 491771 510978 491790
rect 510758 491759 510813 491771
rect 510758 491699 510773 491759
rect 510807 491699 510813 491759
rect 510758 491687 510813 491699
rect 510925 491759 510978 491771
rect 510925 491699 510931 491759
rect 510965 491699 510978 491759
rect 510925 491687 510978 491699
rect 510758 491672 510788 491687
rect 510547 491649 510639 491655
rect 510547 491615 510559 491649
rect 510627 491615 510639 491649
rect 510547 491609 510639 491615
rect 510823 491649 510915 491655
rect 510823 491615 510835 491649
rect 510903 491615 510915 491649
rect 510823 491609 510915 491615
rect 510946 491434 510978 491687
rect 511030 491771 511062 491782
rect 511222 491771 511252 491996
rect 511030 491759 511089 491771
rect 511030 491699 511049 491759
rect 511083 491699 511089 491759
rect 511030 491687 511089 491699
rect 511201 491759 511252 491771
rect 511201 491699 511207 491759
rect 511241 491699 511252 491759
rect 511201 491687 511252 491699
rect 511030 491434 511062 491687
rect 511222 491672 511252 491687
rect 511306 491771 511336 491996
rect 511375 491843 511467 491849
rect 511375 491809 511387 491843
rect 511455 491809 511467 491843
rect 511375 491803 511467 491809
rect 511496 491771 511528 491790
rect 511306 491759 511365 491771
rect 511306 491699 511325 491759
rect 511359 491699 511365 491759
rect 511306 491687 511365 491699
rect 511477 491759 511528 491771
rect 511477 491699 511483 491759
rect 511517 491699 511528 491759
rect 511477 491687 511528 491699
rect 511306 491674 511336 491687
rect 511099 491649 511191 491655
rect 511099 491615 511111 491649
rect 511179 491615 511191 491649
rect 511099 491609 511191 491615
rect 511375 491649 511467 491655
rect 511375 491615 511387 491649
rect 511455 491615 511467 491649
rect 511375 491609 511467 491615
rect 511496 491434 511528 491687
rect 511620 491576 511658 491996
rect 512747 491818 512801 491996
rect 512668 491786 512868 491818
rect 512668 491638 512696 491786
rect 512844 491638 512868 491786
rect 512668 491618 512868 491638
rect 420096 491431 420269 491434
rect 420096 491371 420102 491431
rect 420136 491374 420269 491431
rect 508039 491388 511532 491434
rect 511030 491386 511062 491388
rect 420136 491371 420142 491374
rect 420096 491359 420142 491371
rect 419921 491344 419955 491359
rect 419718 491321 419810 491327
rect 419718 491287 419730 491321
rect 419798 491287 419810 491321
rect 419718 491281 419810 491287
rect 419994 491321 420086 491327
rect 419994 491287 420006 491321
rect 420074 491287 420086 491321
rect 419994 491281 420086 491287
rect 420237 491322 420269 491374
rect 509538 491334 509660 491344
rect 420237 491174 420273 491322
rect 419015 491172 420273 491174
rect 419017 491142 420273 491172
rect 509538 491290 509566 491334
rect 509638 491290 509660 491334
rect 419017 491141 419585 491142
rect 419017 491138 419051 491141
rect 419293 491140 419585 491141
rect 509538 491108 509660 491290
rect 510000 491270 510090 491286
rect 510000 491206 510012 491270
rect 510084 491206 510090 491270
rect 509504 491100 509704 491108
rect 418873 491044 419073 491066
rect 322870 489490 323194 490892
rect 418812 490882 419076 491044
rect 419395 490996 419573 491026
rect 412872 490618 419076 490882
rect 419388 490990 419573 490996
rect 419388 490930 419439 490990
rect 419533 490930 419573 490990
rect 419388 490760 419573 490930
rect 508428 490908 509704 491100
rect 508428 490882 509702 490908
rect 502872 490836 509702 490882
rect 322872 489146 323136 489490
rect 412872 489146 413136 490618
rect 419388 490340 419564 490760
rect 502872 490618 508692 490836
rect 417078 489740 421758 490340
rect 247591 488627 249092 488633
rect 52310 479406 52640 480230
rect 53366 479406 53762 480230
rect 52310 478812 53762 479406
rect 142310 480230 143762 485815
rect 142310 479406 142640 480230
rect 143366 479406 143762 480230
rect 142310 478812 143762 479406
rect 232310 480230 233762 487388
rect 232310 479406 232640 480230
rect 233366 479406 233762 480230
rect 232310 478812 233762 479406
rect 322310 480230 323762 489146
rect 322310 479406 322640 480230
rect 323366 479406 323762 480230
rect 322310 478812 323762 479406
rect 412310 480230 413762 489146
rect 417078 488820 418038 489740
rect 417078 488220 417238 488820
rect 417838 488220 418038 488820
rect 417078 488060 418038 488220
rect 420798 488820 421758 489740
rect 502872 489146 503136 490618
rect 510000 490340 510090 491206
rect 507078 490336 509388 490340
rect 509652 490336 511758 490340
rect 507078 489740 511758 490336
rect 420798 488220 420958 488820
rect 421558 488220 421758 488820
rect 420798 488060 421758 488220
rect 412310 479406 412640 480230
rect 413366 479406 413762 480230
rect 412310 478812 413762 479406
rect 502310 480230 503762 489146
rect 507078 488820 508038 489740
rect 507078 488220 507238 488820
rect 507838 488220 508038 488820
rect 507078 488060 508038 488220
rect 510798 488820 511758 489740
rect 510798 488220 510958 488820
rect 511558 488220 511758 488820
rect 510798 488060 511758 488220
rect 502310 479406 502640 480230
rect 503366 479406 503762 480230
rect 502310 478812 503762 479406
rect 64394 384794 65846 385158
rect 64394 383970 64790 384794
rect 65516 383970 65846 384794
rect 64394 378735 65846 383970
rect 154394 384794 155846 385158
rect 154394 383970 154790 384794
rect 155516 383970 155846 384794
rect 154394 378735 155846 383970
rect 244394 384794 245846 385158
rect 244394 383970 244790 384794
rect 245516 383970 245846 384794
rect 244394 375113 245846 383970
rect 334394 384794 335846 385158
rect 334394 383970 334790 384794
rect 335516 383970 335846 384794
rect 334394 374824 335846 383970
rect 424394 384794 425846 385158
rect 424394 383970 424790 384794
rect 425516 383970 425846 384794
rect 417138 375400 418098 375560
rect 417138 374800 417298 375400
rect 417898 374800 418098 375400
rect 417138 373880 418098 374800
rect 420858 375400 421818 375560
rect 420858 374800 421018 375400
rect 421618 374800 421818 375400
rect 424394 374824 425846 383970
rect 514394 384794 515846 385158
rect 514394 383970 514790 384794
rect 515516 383970 515846 384794
rect 507138 375400 508098 375560
rect 420858 373880 421818 374800
rect 323744 373502 324264 373736
rect 323744 373378 323908 373502
rect 324016 373378 324264 373502
rect 230433 372790 231381 372796
rect 51258 371469 52348 372005
rect 68318 371723 69188 371755
rect 53461 371657 69188 371723
rect 53341 371553 53433 371559
rect 53341 371519 53353 371553
rect 53421 371519 53433 371553
rect 53341 371513 53433 371519
rect 53466 371481 53506 371657
rect 53285 371469 53331 371481
rect 51258 371411 53291 371469
rect 51258 369730 52348 371411
rect 53127 371233 53169 371411
rect 53285 371409 53291 371411
rect 53325 371409 53331 371469
rect 53285 371397 53331 371409
rect 53443 371469 53506 371481
rect 53443 371409 53449 371469
rect 53483 371409 53506 371469
rect 53443 371397 53506 371409
rect 53466 371391 53506 371397
rect 53548 371481 53588 371657
rect 53617 371553 53709 371559
rect 53617 371519 53629 371553
rect 53697 371519 53709 371553
rect 53617 371513 53709 371519
rect 53893 371553 53985 371559
rect 53893 371519 53905 371553
rect 53973 371519 53985 371553
rect 53893 371513 53985 371519
rect 53742 371481 53772 371489
rect 53548 371469 53607 371481
rect 53548 371409 53567 371469
rect 53601 371409 53607 371469
rect 53548 371397 53607 371409
rect 53719 371469 53772 371481
rect 53719 371409 53725 371469
rect 53759 371409 53772 371469
rect 53719 371397 53772 371409
rect 53548 371393 53588 371397
rect 53341 371359 53433 371365
rect 53341 371325 53353 371359
rect 53421 371325 53433 371359
rect 53341 371319 53433 371325
rect 53617 371359 53709 371365
rect 53617 371325 53629 371359
rect 53697 371325 53709 371359
rect 53617 371319 53709 371325
rect 53742 371233 53772 371397
rect 53828 371481 53858 371489
rect 54024 371481 54064 371657
rect 53828 371469 53883 371481
rect 53828 371409 53843 371469
rect 53877 371409 53883 371469
rect 53828 371397 53883 371409
rect 53995 371469 54064 371481
rect 53995 371409 54001 371469
rect 54035 371409 54064 371469
rect 53995 371397 54064 371409
rect 53828 371233 53858 371397
rect 54024 371393 54064 371397
rect 54092 371481 54132 371657
rect 54169 371553 54261 371559
rect 54169 371519 54181 371553
rect 54249 371519 54261 371553
rect 54169 371513 54261 371519
rect 54445 371553 54537 371559
rect 54445 371519 54457 371553
rect 54525 371519 54537 371553
rect 54445 371513 54537 371519
rect 54296 371481 54326 371489
rect 54092 371469 54159 371481
rect 54092 371409 54119 371469
rect 54153 371409 54159 371469
rect 54092 371397 54159 371409
rect 54271 371469 54326 371481
rect 54271 371409 54277 371469
rect 54311 371409 54326 371469
rect 54271 371397 54326 371409
rect 54092 371393 54132 371397
rect 53893 371359 53985 371365
rect 53893 371325 53905 371359
rect 53973 371325 53985 371359
rect 53893 371319 53985 371325
rect 54169 371359 54261 371365
rect 54169 371325 54181 371359
rect 54249 371325 54261 371359
rect 54169 371319 54261 371325
rect 54296 371233 54326 371397
rect 54382 371481 54412 371489
rect 54572 371481 54612 371657
rect 54382 371469 54435 371481
rect 54382 371409 54395 371469
rect 54429 371409 54435 371469
rect 54382 371397 54435 371409
rect 54547 371469 54612 371481
rect 54547 371409 54553 371469
rect 54587 371409 54612 371469
rect 54547 371397 54612 371409
rect 54382 371233 54412 371397
rect 54572 371389 54612 371397
rect 54644 371481 54684 371657
rect 54721 371553 54813 371559
rect 54721 371519 54733 371553
rect 54801 371519 54813 371553
rect 54721 371513 54813 371519
rect 54997 371553 55089 371559
rect 54997 371519 55009 371553
rect 55077 371519 55089 371553
rect 54997 371513 55089 371519
rect 54844 371481 54874 371489
rect 54644 371469 54711 371481
rect 54644 371409 54671 371469
rect 54705 371409 54711 371469
rect 54644 371397 54711 371409
rect 54823 371469 54874 371481
rect 54823 371409 54829 371469
rect 54863 371409 54874 371469
rect 54823 371397 54874 371409
rect 54644 371393 54684 371397
rect 54445 371359 54537 371365
rect 54445 371325 54457 371359
rect 54525 371325 54537 371359
rect 54445 371319 54537 371325
rect 54721 371359 54813 371365
rect 54721 371325 54733 371359
rect 54801 371325 54813 371359
rect 54721 371319 54813 371325
rect 54844 371233 54874 371397
rect 54936 371481 54966 371487
rect 55124 371481 55164 371657
rect 54936 371469 54987 371481
rect 54936 371409 54947 371469
rect 54981 371409 54987 371469
rect 54936 371397 54987 371409
rect 55099 371469 55164 371481
rect 55099 371409 55105 371469
rect 55139 371409 55164 371469
rect 55099 371397 55164 371409
rect 55204 371481 55244 371657
rect 55273 371553 55365 371559
rect 55273 371519 55285 371553
rect 55353 371519 55365 371553
rect 55273 371513 55365 371519
rect 55549 371553 55641 371559
rect 55549 371519 55561 371553
rect 55629 371519 55641 371553
rect 55549 371513 55641 371519
rect 55394 371481 55424 371487
rect 55204 371469 55263 371481
rect 55204 371409 55223 371469
rect 55257 371409 55263 371469
rect 55204 371397 55263 371409
rect 55375 371469 55424 371481
rect 55375 371409 55381 371469
rect 55415 371409 55424 371469
rect 55375 371397 55424 371409
rect 54936 371233 54966 371397
rect 54997 371359 55089 371365
rect 54997 371325 55009 371359
rect 55077 371325 55089 371359
rect 54997 371319 55089 371325
rect 55273 371359 55365 371365
rect 55273 371325 55285 371359
rect 55353 371325 55365 371359
rect 55273 371319 55365 371325
rect 55394 371233 55424 371397
rect 55486 371481 55516 371485
rect 55678 371481 55718 371657
rect 55486 371469 55539 371481
rect 55486 371409 55499 371469
rect 55533 371409 55539 371469
rect 55486 371397 55539 371409
rect 55651 371469 55718 371481
rect 55651 371409 55657 371469
rect 55691 371409 55718 371469
rect 55651 371397 55718 371409
rect 55486 371233 55516 371397
rect 55678 371393 55718 371397
rect 55752 371481 55792 371657
rect 55825 371553 55917 371559
rect 55825 371519 55837 371553
rect 55905 371519 55917 371553
rect 55825 371513 55917 371519
rect 56101 371553 56193 371559
rect 56101 371519 56113 371553
rect 56181 371519 56193 371553
rect 56101 371513 56193 371519
rect 55950 371481 55980 371485
rect 55752 371469 55815 371481
rect 55752 371409 55775 371469
rect 55809 371409 55815 371469
rect 55752 371397 55815 371409
rect 55927 371469 55980 371481
rect 55927 371409 55933 371469
rect 55967 371409 55980 371469
rect 55927 371397 55980 371409
rect 55752 371395 55792 371397
rect 55549 371359 55641 371365
rect 55549 371325 55561 371359
rect 55629 371325 55641 371359
rect 55549 371319 55641 371325
rect 55825 371359 55917 371365
rect 55825 371325 55837 371359
rect 55905 371325 55917 371359
rect 55825 371319 55917 371325
rect 55950 371233 55980 371397
rect 56038 371481 56068 371483
rect 56230 371481 56270 371657
rect 56038 371469 56091 371481
rect 56038 371409 56051 371469
rect 56085 371409 56091 371469
rect 56038 371397 56091 371409
rect 56203 371469 56270 371481
rect 56203 371409 56209 371469
rect 56243 371409 56270 371469
rect 56203 371397 56270 371409
rect 56038 371233 56068 371397
rect 56230 371391 56270 371397
rect 56300 371481 56340 371657
rect 56377 371553 56469 371559
rect 56377 371519 56389 371553
rect 56457 371519 56469 371553
rect 56377 371513 56469 371519
rect 56653 371553 56745 371559
rect 56653 371519 56665 371553
rect 56733 371519 56745 371553
rect 56653 371513 56745 371519
rect 56500 371481 56530 371483
rect 56300 371469 56367 371481
rect 56300 371409 56327 371469
rect 56361 371409 56367 371469
rect 56300 371397 56367 371409
rect 56479 371469 56530 371481
rect 56479 371409 56485 371469
rect 56519 371409 56530 371469
rect 56479 371397 56530 371409
rect 56300 371395 56340 371397
rect 56101 371359 56193 371365
rect 56377 371363 56469 371365
rect 56101 371325 56113 371359
rect 56181 371325 56193 371359
rect 56374 371359 56469 371363
rect 56374 371330 56389 371359
rect 56101 371319 56193 371325
rect 56377 371325 56389 371330
rect 56457 371325 56469 371359
rect 56377 371319 56469 371325
rect 56500 371233 56530 371397
rect 56588 371481 56618 371483
rect 56778 371481 56818 371657
rect 56588 371469 56643 371481
rect 56588 371409 56603 371469
rect 56637 371409 56643 371469
rect 56588 371397 56643 371409
rect 56755 371469 56818 371481
rect 56755 371409 56761 371469
rect 56795 371409 56818 371469
rect 56755 371397 56818 371409
rect 56588 371233 56618 371397
rect 56778 371391 56818 371397
rect 56856 371481 56896 371657
rect 56929 371553 57021 371559
rect 56929 371519 56941 371553
rect 57009 371519 57021 371553
rect 56929 371513 57021 371519
rect 57205 371553 57297 371559
rect 57205 371519 57217 371553
rect 57285 371519 57297 371553
rect 57205 371513 57297 371519
rect 57052 371481 57082 371485
rect 56856 371469 56919 371481
rect 56856 371409 56879 371469
rect 56913 371409 56919 371469
rect 56856 371397 56919 371409
rect 57031 371469 57082 371481
rect 57031 371409 57037 371469
rect 57071 371409 57082 371469
rect 57031 371397 57082 371409
rect 56856 371395 56896 371397
rect 56653 371359 56745 371365
rect 56653 371325 56665 371359
rect 56733 371325 56745 371359
rect 56653 371319 56745 371325
rect 56929 371359 57021 371365
rect 56929 371325 56941 371359
rect 57009 371325 57021 371359
rect 56929 371319 57021 371325
rect 57052 371233 57082 371397
rect 57140 371481 57170 371485
rect 57332 371481 57372 371657
rect 57140 371469 57195 371481
rect 57140 371409 57155 371469
rect 57189 371409 57195 371469
rect 57140 371397 57195 371409
rect 57307 371469 57372 371481
rect 57307 371409 57313 371469
rect 57347 371409 57372 371469
rect 57307 371397 57372 371409
rect 57140 371233 57170 371397
rect 57332 371383 57372 371397
rect 57410 371481 57450 371657
rect 57481 371553 57573 371559
rect 57481 371519 57493 371553
rect 57561 371519 57573 371553
rect 57481 371513 57573 371519
rect 57757 371553 57849 371559
rect 57757 371519 57769 371553
rect 57837 371519 57849 371553
rect 57757 371513 57849 371519
rect 57604 371481 57634 371485
rect 57410 371469 57471 371481
rect 57410 371409 57431 371469
rect 57465 371409 57471 371469
rect 57410 371397 57471 371409
rect 57583 371469 57634 371481
rect 57583 371409 57589 371469
rect 57623 371409 57634 371469
rect 57583 371397 57634 371409
rect 57410 371391 57450 371397
rect 57205 371359 57297 371365
rect 57205 371325 57217 371359
rect 57285 371325 57297 371359
rect 57205 371319 57297 371325
rect 57481 371359 57573 371365
rect 57481 371325 57493 371359
rect 57561 371325 57573 371359
rect 57481 371319 57573 371325
rect 57604 371233 57634 371397
rect 57696 371481 57726 371485
rect 57888 371481 57928 371657
rect 57696 371469 57747 371481
rect 57696 371409 57707 371469
rect 57741 371409 57747 371469
rect 57696 371397 57747 371409
rect 57859 371469 57928 371481
rect 57859 371409 57865 371469
rect 57899 371409 57928 371469
rect 57859 371397 57928 371409
rect 57962 371481 58002 371657
rect 58033 371553 58125 371559
rect 58033 371519 58045 371553
rect 58113 371519 58125 371553
rect 58033 371513 58125 371519
rect 58309 371553 58401 371559
rect 58309 371519 58321 371553
rect 58389 371519 58401 371553
rect 58309 371513 58401 371519
rect 58158 371481 58188 371495
rect 57962 371469 58023 371481
rect 57962 371409 57983 371469
rect 58017 371409 58023 371469
rect 57962 371397 58023 371409
rect 58135 371469 58188 371481
rect 58135 371409 58141 371469
rect 58175 371409 58188 371469
rect 58135 371397 58188 371409
rect 57696 371233 57726 371397
rect 57888 371393 57928 371397
rect 57757 371359 57849 371365
rect 57757 371325 57769 371359
rect 57837 371325 57849 371359
rect 57757 371319 57849 371325
rect 58033 371359 58125 371365
rect 58033 371325 58045 371359
rect 58113 371325 58125 371359
rect 58033 371319 58125 371325
rect 58158 371233 58188 371397
rect 58244 371481 58274 371493
rect 58432 371481 58466 371657
rect 58244 371469 58299 371481
rect 58244 371409 58259 371469
rect 58293 371409 58299 371469
rect 58244 371397 58299 371409
rect 58411 371469 58466 371481
rect 58411 371409 58417 371469
rect 58451 371409 58466 371469
rect 58411 371397 58466 371409
rect 58244 371233 58274 371397
rect 58432 371393 58466 371397
rect 58522 371481 58556 371657
rect 58585 371553 58677 371559
rect 58585 371519 58597 371553
rect 58665 371519 58677 371553
rect 58585 371513 58677 371519
rect 58861 371553 58953 371559
rect 58861 371519 58873 371553
rect 58941 371519 58953 371553
rect 58861 371513 58953 371519
rect 58712 371481 58742 371491
rect 58522 371469 58575 371481
rect 58522 371409 58535 371469
rect 58569 371409 58575 371469
rect 58522 371397 58575 371409
rect 58687 371469 58742 371481
rect 58687 371409 58693 371469
rect 58727 371409 58742 371469
rect 58687 371397 58742 371409
rect 58522 371393 58556 371397
rect 58309 371359 58401 371365
rect 58309 371325 58321 371359
rect 58389 371325 58401 371359
rect 58309 371319 58401 371325
rect 58585 371359 58677 371365
rect 58585 371325 58597 371359
rect 58665 371325 58677 371359
rect 58585 371319 58677 371325
rect 58712 371233 58742 371397
rect 58798 371481 58828 371491
rect 58988 371481 59022 371657
rect 58798 371469 58851 371481
rect 58798 371409 58811 371469
rect 58845 371409 58851 371469
rect 58798 371397 58851 371409
rect 58963 371469 59022 371481
rect 58963 371409 58969 371469
rect 59003 371409 59022 371469
rect 58963 371397 59022 371409
rect 59072 371481 59106 371657
rect 59137 371553 59229 371559
rect 59137 371519 59149 371553
rect 59217 371519 59229 371553
rect 59137 371513 59229 371519
rect 59264 371481 59298 371495
rect 59072 371469 59127 371481
rect 59072 371409 59087 371469
rect 59121 371409 59127 371469
rect 59072 371397 59127 371409
rect 59239 371469 59298 371481
rect 59239 371409 59245 371469
rect 59279 371409 59298 371469
rect 59239 371397 59298 371409
rect 58798 371233 58828 371397
rect 58988 371393 59022 371397
rect 58861 371359 58953 371365
rect 58861 371325 58873 371359
rect 58941 371325 58953 371359
rect 58861 371319 58953 371325
rect 59137 371359 59229 371365
rect 59137 371325 59149 371359
rect 59217 371325 59229 371359
rect 59137 371319 59229 371325
rect 59264 371233 59298 371397
rect 59346 371481 59380 371657
rect 59413 371553 59505 371559
rect 59413 371519 59425 371553
rect 59493 371519 59505 371553
rect 59413 371513 59505 371519
rect 59689 371553 59781 371559
rect 59689 371519 59701 371553
rect 59769 371519 59781 371553
rect 59689 371513 59781 371519
rect 59538 371481 59568 371493
rect 59346 371469 59403 371481
rect 59346 371409 59363 371469
rect 59397 371409 59403 371469
rect 59346 371397 59403 371409
rect 59515 371469 59568 371481
rect 59515 371409 59521 371469
rect 59555 371409 59568 371469
rect 59515 371397 59568 371409
rect 59346 371395 59380 371397
rect 59413 371359 59505 371365
rect 59413 371325 59425 371359
rect 59493 371325 59505 371359
rect 59413 371319 59505 371325
rect 59538 371233 59568 371397
rect 59626 371481 59656 371495
rect 59816 371481 59850 371657
rect 59626 371469 59679 371481
rect 59626 371409 59639 371469
rect 59673 371409 59679 371469
rect 59626 371397 59679 371409
rect 59791 371469 59850 371481
rect 59791 371409 59797 371469
rect 59831 371409 59850 371469
rect 59791 371397 59850 371409
rect 59902 371481 59936 371657
rect 59974 371595 60189 371605
rect 59974 371559 60104 371595
rect 59965 371553 60104 371559
rect 59965 371519 59977 371553
rect 60045 371535 60104 371553
rect 60164 371535 60189 371595
rect 60045 371525 60189 371535
rect 60241 371553 60333 371559
rect 60045 371519 60057 371525
rect 59965 371513 60057 371519
rect 60241 371519 60253 371553
rect 60321 371519 60333 371553
rect 60241 371513 60333 371519
rect 60086 371481 60116 371495
rect 59902 371469 59955 371481
rect 59902 371409 59915 371469
rect 59949 371409 59955 371469
rect 59902 371397 59955 371409
rect 60067 371469 60116 371481
rect 60067 371409 60073 371469
rect 60107 371409 60116 371469
rect 60067 371397 60116 371409
rect 59626 371233 59656 371397
rect 59902 371391 59936 371397
rect 59689 371359 59781 371365
rect 59689 371325 59701 371359
rect 59769 371325 59781 371359
rect 59965 371359 60057 371365
rect 59965 371340 59977 371359
rect 59689 371319 59781 371325
rect 59829 371335 59977 371340
rect 59829 371280 59839 371335
rect 59904 371325 59977 371335
rect 60045 371325 60057 371359
rect 59904 371319 60057 371325
rect 59904 371290 60044 371319
rect 59904 371280 59914 371290
rect 59829 371275 59914 371280
rect 60086 371233 60116 371397
rect 60178 371481 60208 371495
rect 60368 371481 60402 371657
rect 60178 371469 60231 371481
rect 60178 371409 60191 371469
rect 60225 371409 60231 371469
rect 60178 371397 60231 371409
rect 60343 371469 60402 371481
rect 60343 371409 60349 371469
rect 60383 371409 60402 371469
rect 60343 371399 60402 371409
rect 60454 371481 60488 371657
rect 60517 371553 60609 371559
rect 60517 371519 60529 371553
rect 60597 371519 60609 371553
rect 60517 371513 60609 371519
rect 60793 371553 60885 371559
rect 60793 371519 60805 371553
rect 60873 371519 60885 371553
rect 60793 371513 60885 371519
rect 60640 371481 60670 371495
rect 60454 371469 60507 371481
rect 60454 371409 60467 371469
rect 60501 371409 60507 371469
rect 60343 371397 60389 371399
rect 60454 371397 60507 371409
rect 60619 371469 60670 371481
rect 60619 371409 60625 371469
rect 60659 371409 60670 371469
rect 60619 371397 60670 371409
rect 60178 371233 60208 371397
rect 60454 371395 60488 371397
rect 60241 371359 60333 371365
rect 60241 371325 60253 371359
rect 60321 371325 60333 371359
rect 60241 371319 60333 371325
rect 60517 371359 60609 371365
rect 60517 371325 60529 371359
rect 60597 371325 60609 371359
rect 60517 371319 60609 371325
rect 60640 371233 60670 371397
rect 60732 371481 60762 371495
rect 60918 371481 60952 371657
rect 60732 371469 60783 371481
rect 60732 371409 60743 371469
rect 60777 371409 60783 371469
rect 60732 371397 60783 371409
rect 60895 371469 60952 371481
rect 60895 371409 60901 371469
rect 60935 371409 60952 371469
rect 60895 371397 60952 371409
rect 60732 371233 60762 371397
rect 60918 371395 60952 371397
rect 61006 371481 61040 371657
rect 61069 371553 61161 371559
rect 61069 371519 61081 371553
rect 61149 371519 61161 371553
rect 61069 371513 61161 371519
rect 61345 371553 61437 371559
rect 61345 371519 61357 371553
rect 61425 371519 61437 371553
rect 61345 371513 61437 371519
rect 61192 371481 61222 371495
rect 61006 371469 61059 371481
rect 61006 371409 61019 371469
rect 61053 371409 61059 371469
rect 61006 371397 61059 371409
rect 61171 371469 61222 371481
rect 61171 371409 61177 371469
rect 61211 371409 61222 371469
rect 61171 371397 61222 371409
rect 61006 371393 61040 371397
rect 60793 371359 60885 371365
rect 60793 371325 60805 371359
rect 60873 371325 60885 371359
rect 60793 371319 60885 371325
rect 61069 371359 61161 371365
rect 61069 371325 61081 371359
rect 61149 371325 61161 371359
rect 61069 371319 61161 371325
rect 61192 371233 61222 371397
rect 61278 371481 61308 371495
rect 61474 371481 61508 371657
rect 61278 371469 61335 371481
rect 61278 371409 61295 371469
rect 61329 371409 61335 371469
rect 61278 371397 61335 371409
rect 61447 371469 61508 371481
rect 61447 371409 61453 371469
rect 61487 371409 61508 371469
rect 61447 371397 61508 371409
rect 61278 371233 61308 371397
rect 61474 371389 61508 371397
rect 61556 371481 61590 371657
rect 61621 371553 61713 371559
rect 61621 371519 61633 371553
rect 61701 371519 61713 371553
rect 61621 371513 61713 371519
rect 61897 371553 61989 371559
rect 61897 371519 61909 371553
rect 61977 371519 61989 371553
rect 61897 371513 61989 371519
rect 61746 371481 61776 371495
rect 61556 371469 61611 371481
rect 61556 371409 61571 371469
rect 61605 371409 61611 371469
rect 61556 371397 61611 371409
rect 61723 371469 61776 371481
rect 61723 371409 61729 371469
rect 61763 371409 61776 371469
rect 61723 371397 61776 371409
rect 61556 371395 61590 371397
rect 61345 371359 61437 371365
rect 61345 371325 61357 371359
rect 61425 371325 61437 371359
rect 61345 371319 61437 371325
rect 61621 371359 61713 371365
rect 61621 371325 61633 371359
rect 61701 371325 61713 371359
rect 61621 371319 61713 371325
rect 61746 371233 61776 371397
rect 61834 371481 61864 371493
rect 62028 371481 62062 371657
rect 61834 371469 61887 371481
rect 61834 371409 61847 371469
rect 61881 371409 61887 371469
rect 61834 371397 61887 371409
rect 61999 371469 62062 371481
rect 61999 371409 62005 371469
rect 62039 371409 62062 371469
rect 61999 371397 62062 371409
rect 61834 371233 61864 371397
rect 62028 371393 62062 371397
rect 62106 371481 62140 371657
rect 62173 371553 62265 371559
rect 62173 371519 62185 371553
rect 62253 371519 62265 371553
rect 62173 371513 62265 371519
rect 62449 371553 62541 371559
rect 62449 371519 62461 371553
rect 62529 371519 62541 371553
rect 62449 371513 62541 371519
rect 62298 371481 62328 371497
rect 62106 371469 62163 371481
rect 62106 371409 62123 371469
rect 62157 371409 62163 371469
rect 62106 371397 62163 371409
rect 62275 371469 62328 371481
rect 62275 371409 62281 371469
rect 62315 371409 62328 371469
rect 62275 371397 62328 371409
rect 62106 371395 62140 371397
rect 61897 371359 61989 371365
rect 61897 371325 61909 371359
rect 61977 371325 61989 371359
rect 61897 371319 61989 371325
rect 62173 371359 62265 371365
rect 62173 371325 62185 371359
rect 62253 371325 62265 371359
rect 62173 371319 62265 371325
rect 62298 371233 62328 371397
rect 62386 371481 62416 371497
rect 62584 371481 62618 371657
rect 62386 371469 62439 371481
rect 62386 371409 62399 371469
rect 62433 371409 62439 371469
rect 62386 371397 62439 371409
rect 62551 371469 62618 371481
rect 62551 371409 62557 371469
rect 62591 371409 62618 371469
rect 62551 371397 62618 371409
rect 62386 371233 62416 371397
rect 62584 371385 62618 371397
rect 62658 371481 62692 371657
rect 62725 371553 62817 371559
rect 62725 371519 62737 371553
rect 62805 371519 62817 371553
rect 62725 371513 62817 371519
rect 63001 371553 63093 371559
rect 63001 371519 63013 371553
rect 63081 371519 63093 371553
rect 63001 371513 63093 371519
rect 62848 371481 62878 371499
rect 62658 371469 62715 371481
rect 62658 371409 62675 371469
rect 62709 371409 62715 371469
rect 62658 371397 62715 371409
rect 62827 371469 62878 371481
rect 62827 371409 62833 371469
rect 62867 371409 62878 371469
rect 62827 371397 62878 371409
rect 62658 371389 62692 371397
rect 62449 371359 62541 371365
rect 62449 371325 62461 371359
rect 62529 371325 62541 371359
rect 62449 371319 62541 371325
rect 62725 371359 62817 371365
rect 62725 371325 62737 371359
rect 62805 371325 62817 371359
rect 62725 371319 62817 371325
rect 62848 371233 62878 371397
rect 62936 371481 62966 371497
rect 63128 371481 63162 371657
rect 62936 371469 62991 371481
rect 62936 371409 62951 371469
rect 62985 371409 62991 371469
rect 62936 371397 62991 371409
rect 63103 371469 63162 371481
rect 63103 371409 63109 371469
rect 63143 371409 63162 371469
rect 63103 371397 63162 371409
rect 62936 371233 62966 371397
rect 63128 371385 63162 371397
rect 63208 371481 63242 371657
rect 63277 371553 63369 371559
rect 63277 371519 63289 371553
rect 63357 371519 63369 371553
rect 63277 371513 63369 371519
rect 63553 371553 63645 371559
rect 63553 371519 63565 371553
rect 63633 371519 63645 371553
rect 63553 371513 63645 371519
rect 63400 371481 63430 371497
rect 63208 371469 63267 371481
rect 63208 371409 63227 371469
rect 63261 371409 63267 371469
rect 63208 371397 63267 371409
rect 63379 371469 63430 371481
rect 63379 371409 63385 371469
rect 63419 371409 63430 371469
rect 63379 371397 63430 371409
rect 63208 371383 63242 371397
rect 63001 371359 63093 371365
rect 63001 371325 63013 371359
rect 63081 371325 63093 371359
rect 63001 371319 63093 371325
rect 63277 371359 63369 371365
rect 63277 371325 63289 371359
rect 63357 371325 63369 371359
rect 63277 371319 63369 371325
rect 63400 371233 63430 371397
rect 63488 371481 63518 371499
rect 63684 371481 63718 371657
rect 63488 371469 63543 371481
rect 63488 371409 63503 371469
rect 63537 371409 63543 371469
rect 63488 371397 63543 371409
rect 63655 371469 63718 371481
rect 63655 371409 63661 371469
rect 63695 371409 63718 371469
rect 63655 371397 63718 371409
rect 63488 371233 63518 371397
rect 63684 371385 63718 371397
rect 63758 371481 63792 371657
rect 63829 371553 63921 371559
rect 63829 371519 63841 371553
rect 63909 371519 63921 371553
rect 63829 371513 63921 371519
rect 64105 371553 64197 371559
rect 64105 371519 64117 371553
rect 64185 371519 64197 371553
rect 64105 371513 64197 371519
rect 63952 371481 63982 371497
rect 63758 371469 63819 371481
rect 63758 371409 63779 371469
rect 63813 371409 63819 371469
rect 63758 371397 63819 371409
rect 63931 371469 63982 371481
rect 63931 371409 63937 371469
rect 63971 371409 63982 371469
rect 63931 371397 63982 371409
rect 63758 371383 63792 371397
rect 63553 371359 63645 371365
rect 63553 371325 63565 371359
rect 63633 371325 63645 371359
rect 63553 371319 63645 371325
rect 63829 371359 63921 371365
rect 63829 371325 63841 371359
rect 63909 371325 63921 371359
rect 63829 371319 63921 371325
rect 63952 371233 63982 371397
rect 64042 371481 64072 371499
rect 64234 371481 64268 371657
rect 64042 371469 64095 371481
rect 64042 371409 64055 371469
rect 64089 371409 64095 371469
rect 64042 371397 64095 371409
rect 64207 371469 64268 371481
rect 64207 371409 64213 371469
rect 64247 371409 64268 371469
rect 64207 371397 64268 371409
rect 64042 371233 64072 371397
rect 64234 371387 64268 371397
rect 64310 371481 64344 371657
rect 64381 371553 64473 371559
rect 64381 371519 64393 371553
rect 64461 371519 64473 371553
rect 64381 371513 64473 371519
rect 64657 371553 64749 371559
rect 64657 371519 64669 371553
rect 64737 371519 64749 371553
rect 64657 371513 64749 371519
rect 64504 371481 64534 371497
rect 64310 371469 64371 371481
rect 64310 371409 64331 371469
rect 64365 371409 64371 371469
rect 64310 371397 64371 371409
rect 64483 371469 64534 371481
rect 64483 371409 64489 371469
rect 64523 371409 64534 371469
rect 64483 371397 64534 371409
rect 64310 371387 64344 371397
rect 64105 371359 64197 371365
rect 64105 371325 64117 371359
rect 64185 371325 64197 371359
rect 64105 371319 64197 371325
rect 64381 371359 64473 371365
rect 64381 371325 64393 371359
rect 64461 371325 64473 371359
rect 64381 371319 64473 371325
rect 64504 371233 64534 371397
rect 64594 371481 64624 371499
rect 64784 371481 64818 371657
rect 64594 371469 64647 371481
rect 64594 371409 64607 371469
rect 64641 371409 64647 371469
rect 64594 371397 64647 371409
rect 64759 371469 64818 371481
rect 64759 371409 64765 371469
rect 64799 371409 64818 371469
rect 64759 371397 64818 371409
rect 64594 371233 64624 371397
rect 64784 371391 64818 371397
rect 64866 371481 64900 371657
rect 64933 371553 65025 371559
rect 64933 371519 64945 371553
rect 65013 371519 65025 371553
rect 64933 371513 65025 371519
rect 65209 371553 65301 371559
rect 65209 371519 65221 371553
rect 65289 371519 65301 371553
rect 65209 371513 65301 371519
rect 65058 371481 65088 371503
rect 64866 371469 64923 371481
rect 64866 371409 64883 371469
rect 64917 371409 64923 371469
rect 64866 371397 64923 371409
rect 65035 371469 65088 371481
rect 65035 371409 65041 371469
rect 65075 371409 65088 371469
rect 65035 371397 65088 371409
rect 64866 371389 64900 371397
rect 64657 371359 64749 371365
rect 64657 371325 64669 371359
rect 64737 371325 64749 371359
rect 64657 371319 64749 371325
rect 64933 371359 65025 371365
rect 64933 371325 64945 371359
rect 65013 371325 65025 371359
rect 64933 371319 65025 371325
rect 65058 371233 65088 371397
rect 65148 371481 65178 371505
rect 65336 371481 65370 371657
rect 65148 371469 65199 371481
rect 65148 371409 65159 371469
rect 65193 371409 65199 371469
rect 65148 371397 65199 371409
rect 65311 371469 65370 371481
rect 65311 371409 65317 371469
rect 65351 371409 65370 371469
rect 65311 371397 65370 371409
rect 65414 371481 65448 371657
rect 65485 371553 65577 371559
rect 65485 371519 65497 371553
rect 65565 371519 65577 371553
rect 65485 371513 65577 371519
rect 65761 371553 65853 371559
rect 65761 371519 65773 371553
rect 65841 371519 65853 371553
rect 65761 371513 65853 371519
rect 65612 371481 65642 371505
rect 65414 371469 65475 371481
rect 65414 371409 65435 371469
rect 65469 371409 65475 371469
rect 65414 371397 65475 371409
rect 65587 371469 65642 371481
rect 65587 371409 65593 371469
rect 65627 371409 65642 371469
rect 65587 371397 65642 371409
rect 65148 371233 65178 371397
rect 65336 371395 65370 371397
rect 65209 371359 65301 371365
rect 65209 371325 65221 371359
rect 65289 371325 65301 371359
rect 65209 371319 65301 371325
rect 65485 371359 65577 371365
rect 65485 371325 65497 371359
rect 65565 371325 65577 371359
rect 65485 371319 65577 371325
rect 65612 371233 65642 371397
rect 65698 371481 65728 371509
rect 65886 371481 65920 371657
rect 65698 371469 65751 371481
rect 65698 371409 65711 371469
rect 65745 371409 65751 371469
rect 65698 371397 65751 371409
rect 65863 371469 65920 371481
rect 65863 371409 65869 371469
rect 65903 371409 65920 371469
rect 65863 371397 65920 371409
rect 65698 371233 65728 371397
rect 65886 371393 65920 371397
rect 65970 371481 66004 371657
rect 66037 371553 66129 371559
rect 66037 371519 66049 371553
rect 66117 371519 66129 371553
rect 66037 371513 66129 371519
rect 66313 371553 66405 371559
rect 66313 371519 66325 371553
rect 66393 371519 66405 371553
rect 66313 371513 66405 371519
rect 66158 371481 66188 371495
rect 65970 371469 66027 371481
rect 65970 371409 65987 371469
rect 66021 371409 66027 371469
rect 65970 371397 66027 371409
rect 66139 371469 66188 371481
rect 66139 371409 66145 371469
rect 66179 371409 66188 371469
rect 66139 371397 66188 371409
rect 65970 371391 66004 371397
rect 65761 371359 65853 371365
rect 65761 371325 65773 371359
rect 65841 371325 65853 371359
rect 65761 371319 65853 371325
rect 66037 371359 66129 371365
rect 66037 371325 66049 371359
rect 66117 371325 66129 371359
rect 66037 371319 66129 371325
rect 66158 371233 66188 371397
rect 66250 371481 66280 371493
rect 66438 371481 66472 371657
rect 66250 371469 66303 371481
rect 66250 371409 66263 371469
rect 66297 371409 66303 371469
rect 66250 371397 66303 371409
rect 66415 371469 66472 371481
rect 66415 371409 66421 371469
rect 66455 371409 66472 371469
rect 66415 371397 66472 371409
rect 66250 371233 66280 371397
rect 66438 371393 66472 371397
rect 66522 371481 66556 371657
rect 66589 371553 66681 371559
rect 66589 371519 66601 371553
rect 66669 371519 66681 371553
rect 66589 371513 66681 371519
rect 66865 371553 66957 371559
rect 66865 371519 66877 371553
rect 66945 371519 66957 371553
rect 66865 371513 66957 371519
rect 66714 371481 66744 371495
rect 66522 371469 66579 371481
rect 66522 371409 66539 371469
rect 66573 371409 66579 371469
rect 66522 371397 66579 371409
rect 66691 371469 66744 371481
rect 66691 371409 66697 371469
rect 66731 371409 66744 371469
rect 66691 371397 66744 371409
rect 66522 371395 66556 371397
rect 66313 371359 66405 371365
rect 66313 371325 66325 371359
rect 66393 371325 66405 371359
rect 66313 371319 66405 371325
rect 66589 371359 66681 371365
rect 66589 371325 66601 371359
rect 66669 371325 66681 371359
rect 66589 371319 66681 371325
rect 66714 371233 66744 371397
rect 66798 371481 66828 371495
rect 66992 371481 67026 371657
rect 66798 371469 66855 371481
rect 66798 371409 66815 371469
rect 66849 371409 66855 371469
rect 66798 371397 66855 371409
rect 66967 371469 67026 371481
rect 66967 371409 66973 371469
rect 67007 371409 67026 371469
rect 66967 371399 67026 371409
rect 67070 371481 67104 371657
rect 67141 371553 67233 371559
rect 67141 371519 67153 371553
rect 67221 371519 67233 371553
rect 67141 371513 67233 371519
rect 67264 371481 67294 371495
rect 67070 371469 67131 371481
rect 67070 371409 67091 371469
rect 67125 371409 67131 371469
rect 66967 371397 67013 371399
rect 67070 371397 67131 371409
rect 67243 371469 67294 371481
rect 67243 371409 67249 371469
rect 67283 371409 67294 371469
rect 67243 371397 67294 371409
rect 67384 371405 67418 371657
rect 66798 371233 66828 371397
rect 66865 371359 66957 371365
rect 66865 371325 66877 371359
rect 66945 371325 66957 371359
rect 66865 371319 66957 371325
rect 67141 371359 67233 371365
rect 67141 371325 67153 371359
rect 67221 371325 67233 371359
rect 67141 371319 67233 371325
rect 67264 371233 67294 371397
rect 53127 371191 67296 371233
rect 67254 371189 67296 371191
rect 57306 371085 57446 371097
rect 57306 371029 57346 371085
rect 57424 371029 57446 371085
rect 57306 370415 57446 371029
rect 68318 370600 69188 371657
rect 51258 368634 52348 368640
rect 53138 370215 57492 370415
rect 53138 365815 53338 370215
rect 68318 369724 69188 369730
rect 141258 371469 142348 372005
rect 323744 372700 324264 373378
rect 417138 373280 421818 373880
rect 507138 374800 507298 375400
rect 507898 374800 508098 375400
rect 507138 373880 508098 374800
rect 510858 375400 511818 375560
rect 510858 374800 511018 375400
rect 511618 374800 511818 375400
rect 514394 374824 515846 383970
rect 510858 373880 511818 374800
rect 507138 373280 511818 373880
rect 323888 372598 323972 372700
rect 419380 372678 419564 373280
rect 323888 372556 323904 372598
rect 323958 372556 323972 372598
rect 419368 372592 420088 372678
rect 323888 372536 323972 372556
rect 338790 372400 339590 372534
rect 321787 372028 321793 372354
rect 322119 372146 322656 372354
rect 324001 372334 339590 372400
rect 323881 372231 323973 372237
rect 323881 372197 323893 372231
rect 323961 372197 323973 372231
rect 323881 372191 323973 372197
rect 324006 372159 324046 372334
rect 323825 372147 323871 372159
rect 323825 372146 323831 372147
rect 322119 372088 323831 372146
rect 322119 372028 322656 372088
rect 323667 371910 323709 372088
rect 323825 372087 323831 372088
rect 323865 372087 323871 372147
rect 323825 372075 323871 372087
rect 323983 372147 324046 372159
rect 323983 372087 323989 372147
rect 324023 372087 324046 372147
rect 323983 372075 324046 372087
rect 324006 372068 324046 372075
rect 324088 372159 324128 372334
rect 324157 372231 324249 372237
rect 324157 372197 324169 372231
rect 324237 372197 324249 372231
rect 324157 372191 324249 372197
rect 324433 372231 324525 372237
rect 324433 372197 324445 372231
rect 324513 372197 324525 372231
rect 324433 372191 324525 372197
rect 324282 372159 324312 372166
rect 324088 372147 324147 372159
rect 324088 372087 324107 372147
rect 324141 372087 324147 372147
rect 324088 372075 324147 372087
rect 324259 372147 324312 372159
rect 324259 372087 324265 372147
rect 324299 372087 324312 372147
rect 324259 372075 324312 372087
rect 324088 372070 324128 372075
rect 323881 372037 323973 372043
rect 323881 372003 323893 372037
rect 323961 372003 323973 372037
rect 323881 371997 323973 372003
rect 324157 372037 324249 372043
rect 324157 372003 324169 372037
rect 324237 372003 324249 372037
rect 324157 371997 324249 372003
rect 323839 371910 324015 371911
rect 324282 371910 324312 372075
rect 324368 372159 324398 372166
rect 324564 372159 324604 372334
rect 324368 372147 324423 372159
rect 324368 372087 324383 372147
rect 324417 372087 324423 372147
rect 324368 372075 324423 372087
rect 324535 372147 324604 372159
rect 324535 372087 324541 372147
rect 324575 372087 324604 372147
rect 324535 372075 324604 372087
rect 324368 371910 324398 372075
rect 324564 372070 324604 372075
rect 324632 372159 324672 372334
rect 324709 372231 324801 372237
rect 324709 372197 324721 372231
rect 324789 372197 324801 372231
rect 324709 372191 324801 372197
rect 324985 372231 325077 372237
rect 324985 372197 324997 372231
rect 325065 372197 325077 372231
rect 324985 372191 325077 372197
rect 324836 372159 324866 372166
rect 324632 372147 324699 372159
rect 324632 372087 324659 372147
rect 324693 372087 324699 372147
rect 324632 372075 324699 372087
rect 324811 372147 324866 372159
rect 324811 372087 324817 372147
rect 324851 372087 324866 372147
rect 324811 372075 324866 372087
rect 324632 372070 324672 372075
rect 324433 372037 324525 372043
rect 324433 372003 324445 372037
rect 324513 372003 324525 372037
rect 324433 371997 324525 372003
rect 324709 372037 324801 372043
rect 324709 372003 324721 372037
rect 324789 372003 324801 372037
rect 324709 371997 324801 372003
rect 324836 371910 324866 372075
rect 324922 372159 324952 372166
rect 325112 372159 325152 372334
rect 324922 372147 324975 372159
rect 324922 372087 324935 372147
rect 324969 372087 324975 372147
rect 324922 372075 324975 372087
rect 325087 372147 325152 372159
rect 325087 372087 325093 372147
rect 325127 372087 325152 372147
rect 325087 372075 325152 372087
rect 324922 371910 324952 372075
rect 325112 372066 325152 372075
rect 325184 372159 325224 372334
rect 325261 372231 325353 372237
rect 325261 372197 325273 372231
rect 325341 372197 325353 372231
rect 325261 372191 325353 372197
rect 325537 372231 325629 372237
rect 325537 372197 325549 372231
rect 325617 372197 325629 372231
rect 325537 372191 325629 372197
rect 325384 372159 325414 372166
rect 325184 372147 325251 372159
rect 325184 372087 325211 372147
rect 325245 372087 325251 372147
rect 325184 372075 325251 372087
rect 325363 372147 325414 372159
rect 325363 372087 325369 372147
rect 325403 372087 325414 372147
rect 325363 372075 325414 372087
rect 325184 372070 325224 372075
rect 324985 372037 325077 372043
rect 324985 372003 324997 372037
rect 325065 372003 325077 372037
rect 324985 371997 325077 372003
rect 325261 372037 325353 372043
rect 325261 372003 325273 372037
rect 325341 372003 325353 372037
rect 325261 371997 325353 372003
rect 325384 371910 325414 372075
rect 325476 372159 325506 372164
rect 325664 372159 325704 372334
rect 325476 372147 325527 372159
rect 325476 372087 325487 372147
rect 325521 372087 325527 372147
rect 325476 372075 325527 372087
rect 325639 372147 325704 372159
rect 325639 372087 325645 372147
rect 325679 372087 325704 372147
rect 325639 372075 325704 372087
rect 325476 371910 325506 372075
rect 325664 372074 325704 372075
rect 325744 372159 325784 372334
rect 325813 372231 325905 372237
rect 325813 372197 325825 372231
rect 325893 372197 325905 372231
rect 325813 372191 325905 372197
rect 326089 372231 326181 372237
rect 326089 372197 326101 372231
rect 326169 372197 326181 372231
rect 326089 372191 326181 372197
rect 325934 372159 325964 372164
rect 325744 372147 325803 372159
rect 325744 372087 325763 372147
rect 325797 372087 325803 372147
rect 325744 372075 325803 372087
rect 325915 372147 325964 372159
rect 325915 372087 325921 372147
rect 325955 372087 325964 372147
rect 325915 372075 325964 372087
rect 325744 372074 325784 372075
rect 325537 372037 325629 372043
rect 325537 372003 325549 372037
rect 325617 372003 325629 372037
rect 325537 371997 325629 372003
rect 325813 372037 325905 372043
rect 325813 372003 325825 372037
rect 325893 372003 325905 372037
rect 325813 371997 325905 372003
rect 325934 371910 325964 372075
rect 326026 372159 326056 372162
rect 326218 372159 326258 372334
rect 326026 372147 326079 372159
rect 326026 372087 326039 372147
rect 326073 372087 326079 372147
rect 326026 372075 326079 372087
rect 326191 372147 326258 372159
rect 326191 372087 326197 372147
rect 326231 372087 326258 372147
rect 326191 372075 326258 372087
rect 326026 371910 326056 372075
rect 326218 372070 326258 372075
rect 326292 372159 326332 372334
rect 326365 372231 326457 372237
rect 326365 372197 326377 372231
rect 326445 372197 326457 372231
rect 326365 372191 326457 372197
rect 326641 372231 326733 372237
rect 326641 372197 326653 372231
rect 326721 372197 326733 372231
rect 326641 372191 326733 372197
rect 326490 372159 326520 372162
rect 326292 372147 326355 372159
rect 326292 372087 326315 372147
rect 326349 372087 326355 372147
rect 326292 372075 326355 372087
rect 326467 372147 326520 372159
rect 326467 372087 326473 372147
rect 326507 372087 326520 372147
rect 326467 372075 326520 372087
rect 326292 372072 326332 372075
rect 326089 372037 326181 372043
rect 326089 372003 326101 372037
rect 326169 372003 326181 372037
rect 326089 371997 326181 372003
rect 326365 372037 326457 372043
rect 326365 372003 326377 372037
rect 326445 372003 326457 372037
rect 326365 371997 326457 372003
rect 326490 371910 326520 372075
rect 326578 372159 326608 372160
rect 326770 372159 326810 372334
rect 326578 372147 326631 372159
rect 326578 372087 326591 372147
rect 326625 372087 326631 372147
rect 326578 372075 326631 372087
rect 326743 372147 326810 372159
rect 326743 372087 326749 372147
rect 326783 372087 326810 372147
rect 326743 372075 326810 372087
rect 326578 371910 326608 372075
rect 326770 372068 326810 372075
rect 326840 372159 326880 372334
rect 326917 372231 327009 372237
rect 326917 372197 326929 372231
rect 326997 372197 327009 372231
rect 326917 372191 327009 372197
rect 327193 372231 327285 372237
rect 327193 372197 327205 372231
rect 327273 372197 327285 372231
rect 327193 372191 327285 372197
rect 327040 372159 327070 372160
rect 326840 372147 326907 372159
rect 326840 372087 326867 372147
rect 326901 372087 326907 372147
rect 326840 372075 326907 372087
rect 327019 372147 327070 372159
rect 327019 372087 327025 372147
rect 327059 372087 327070 372147
rect 327019 372075 327070 372087
rect 326840 372072 326880 372075
rect 326641 372037 326733 372043
rect 326641 372003 326653 372037
rect 326721 372003 326733 372037
rect 326641 371997 326733 372003
rect 326917 372037 327009 372043
rect 326917 372003 326929 372037
rect 326997 372003 327009 372037
rect 326917 371997 327009 372003
rect 327040 371910 327070 372075
rect 327128 372159 327158 372160
rect 327318 372159 327358 372334
rect 327128 372147 327183 372159
rect 327128 372087 327143 372147
rect 327177 372087 327183 372147
rect 327128 372075 327183 372087
rect 327295 372147 327358 372159
rect 327295 372087 327301 372147
rect 327335 372087 327358 372147
rect 327295 372075 327358 372087
rect 327128 371910 327158 372075
rect 327318 372068 327358 372075
rect 327396 372159 327436 372334
rect 327469 372231 327561 372237
rect 327469 372197 327481 372231
rect 327549 372197 327561 372231
rect 327469 372191 327561 372197
rect 327745 372231 327837 372237
rect 327745 372197 327757 372231
rect 327825 372197 327837 372231
rect 327745 372191 327837 372197
rect 327592 372159 327622 372162
rect 327396 372147 327459 372159
rect 327396 372087 327419 372147
rect 327453 372087 327459 372147
rect 327396 372075 327459 372087
rect 327571 372147 327622 372159
rect 327571 372087 327577 372147
rect 327611 372087 327622 372147
rect 327571 372075 327622 372087
rect 327396 372072 327436 372075
rect 327193 372037 327285 372043
rect 327193 372003 327205 372037
rect 327273 372003 327285 372037
rect 327193 371997 327285 372003
rect 327469 372037 327561 372043
rect 327469 372003 327481 372037
rect 327549 372003 327561 372037
rect 327469 371997 327561 372003
rect 327592 371910 327622 372075
rect 327680 372159 327710 372162
rect 327872 372159 327912 372334
rect 327680 372147 327735 372159
rect 327680 372087 327695 372147
rect 327729 372087 327735 372147
rect 327680 372075 327735 372087
rect 327847 372147 327912 372159
rect 327847 372087 327853 372147
rect 327887 372087 327912 372147
rect 327847 372075 327912 372087
rect 327680 371910 327710 372075
rect 327872 372060 327912 372075
rect 327950 372159 327990 372334
rect 328021 372231 328113 372237
rect 328021 372197 328033 372231
rect 328101 372197 328113 372231
rect 328021 372191 328113 372197
rect 328297 372231 328389 372237
rect 328297 372197 328309 372231
rect 328377 372197 328389 372231
rect 328297 372191 328389 372197
rect 328144 372159 328174 372162
rect 327950 372147 328011 372159
rect 327950 372087 327971 372147
rect 328005 372087 328011 372147
rect 327950 372075 328011 372087
rect 328123 372147 328174 372159
rect 328123 372087 328129 372147
rect 328163 372087 328174 372147
rect 328123 372075 328174 372087
rect 327950 372068 327990 372075
rect 327745 372037 327837 372043
rect 327745 372003 327757 372037
rect 327825 372003 327837 372037
rect 327745 371997 327837 372003
rect 328021 372037 328113 372043
rect 328021 372003 328033 372037
rect 328101 372003 328113 372037
rect 328021 371997 328113 372003
rect 328144 371910 328174 372075
rect 328236 372159 328266 372162
rect 328428 372159 328468 372334
rect 328236 372147 328287 372159
rect 328236 372087 328247 372147
rect 328281 372087 328287 372147
rect 328236 372075 328287 372087
rect 328399 372147 328468 372159
rect 328399 372087 328405 372147
rect 328439 372087 328468 372147
rect 328399 372075 328468 372087
rect 328236 371910 328266 372075
rect 328428 372070 328468 372075
rect 328502 372159 328542 372334
rect 328573 372231 328665 372237
rect 328573 372197 328585 372231
rect 328653 372197 328665 372231
rect 328573 372191 328665 372197
rect 328849 372231 328941 372237
rect 328849 372197 328861 372231
rect 328929 372197 328941 372231
rect 328849 372191 328941 372197
rect 328698 372159 328728 372172
rect 328502 372147 328563 372159
rect 328502 372087 328523 372147
rect 328557 372087 328563 372147
rect 328502 372075 328563 372087
rect 328675 372147 328728 372159
rect 328675 372087 328681 372147
rect 328715 372087 328728 372147
rect 328675 372075 328728 372087
rect 328502 372074 328542 372075
rect 328297 372037 328389 372043
rect 328297 372003 328309 372037
rect 328377 372003 328389 372037
rect 328297 371997 328389 372003
rect 328573 372037 328665 372043
rect 328573 372003 328585 372037
rect 328653 372003 328665 372037
rect 328573 371997 328665 372003
rect 328698 371910 328728 372075
rect 328784 372159 328814 372170
rect 328972 372159 329006 372334
rect 328784 372147 328839 372159
rect 328784 372087 328799 372147
rect 328833 372087 328839 372147
rect 328784 372075 328839 372087
rect 328951 372147 329006 372159
rect 328951 372087 328957 372147
rect 328991 372087 329006 372147
rect 328951 372075 329006 372087
rect 328784 371910 328814 372075
rect 328972 372070 329006 372075
rect 329062 372159 329096 372334
rect 329125 372231 329217 372237
rect 329125 372197 329137 372231
rect 329205 372197 329217 372231
rect 329125 372191 329217 372197
rect 329401 372231 329493 372237
rect 329401 372197 329413 372231
rect 329481 372197 329493 372231
rect 329401 372191 329493 372197
rect 329252 372159 329282 372168
rect 329062 372147 329115 372159
rect 329062 372087 329075 372147
rect 329109 372087 329115 372147
rect 329062 372075 329115 372087
rect 329227 372147 329282 372159
rect 329227 372087 329233 372147
rect 329267 372087 329282 372147
rect 329227 372075 329282 372087
rect 329062 372070 329096 372075
rect 328849 372037 328941 372043
rect 328849 372003 328861 372037
rect 328929 372003 328941 372037
rect 328849 371997 328941 372003
rect 329125 372037 329217 372043
rect 329125 372003 329137 372037
rect 329205 372003 329217 372037
rect 329125 371997 329217 372003
rect 329252 371910 329282 372075
rect 329338 372159 329368 372168
rect 329528 372159 329562 372334
rect 329338 372147 329391 372159
rect 329338 372087 329351 372147
rect 329385 372087 329391 372147
rect 329338 372075 329391 372087
rect 329503 372147 329562 372159
rect 329503 372087 329509 372147
rect 329543 372087 329562 372147
rect 329503 372075 329562 372087
rect 329338 371910 329368 372075
rect 329528 372070 329562 372075
rect 329612 372159 329646 372334
rect 329677 372231 329769 372237
rect 329677 372197 329689 372231
rect 329757 372197 329769 372231
rect 329677 372191 329769 372197
rect 329804 372159 329838 372172
rect 329612 372147 329667 372159
rect 329612 372087 329627 372147
rect 329661 372087 329667 372147
rect 329612 372075 329667 372087
rect 329779 372147 329838 372159
rect 329779 372087 329785 372147
rect 329819 372087 329838 372147
rect 329779 372075 329838 372087
rect 329612 372074 329646 372075
rect 329401 372037 329493 372043
rect 329401 372003 329413 372037
rect 329481 372003 329493 372037
rect 329401 371997 329493 372003
rect 329677 372037 329769 372043
rect 329677 372003 329689 372037
rect 329757 372003 329769 372037
rect 329677 371997 329769 372003
rect 329804 371910 329838 372075
rect 329886 372159 329920 372334
rect 329953 372231 330045 372237
rect 329953 372197 329965 372231
rect 330033 372197 330045 372231
rect 329953 372191 330045 372197
rect 330229 372231 330321 372237
rect 330229 372197 330241 372231
rect 330309 372197 330321 372231
rect 330229 372191 330321 372197
rect 330078 372159 330108 372170
rect 329886 372147 329943 372159
rect 329886 372087 329903 372147
rect 329937 372087 329943 372147
rect 329886 372075 329943 372087
rect 330055 372147 330108 372159
rect 330055 372087 330061 372147
rect 330095 372087 330108 372147
rect 330055 372075 330108 372087
rect 329886 372072 329920 372075
rect 329953 372037 330045 372043
rect 329953 372003 329965 372037
rect 330033 372003 330045 372037
rect 329953 371997 330045 372003
rect 330078 371910 330108 372075
rect 330166 372159 330196 372172
rect 330356 372159 330390 372334
rect 330166 372147 330219 372159
rect 330166 372087 330179 372147
rect 330213 372087 330219 372147
rect 330166 372075 330219 372087
rect 330331 372147 330390 372159
rect 330331 372087 330337 372147
rect 330371 372087 330390 372147
rect 330331 372075 330390 372087
rect 330166 371910 330196 372075
rect 330356 372074 330390 372075
rect 330442 372159 330476 372334
rect 330505 372231 330597 372237
rect 330505 372197 330517 372231
rect 330585 372197 330597 372231
rect 330505 372191 330597 372197
rect 330781 372231 330873 372237
rect 330781 372197 330793 372231
rect 330861 372197 330873 372231
rect 330781 372191 330873 372197
rect 330626 372159 330656 372172
rect 330442 372147 330495 372159
rect 330442 372087 330455 372147
rect 330489 372087 330495 372147
rect 330442 372075 330495 372087
rect 330607 372147 330656 372159
rect 330607 372087 330613 372147
rect 330647 372087 330656 372147
rect 330607 372075 330656 372087
rect 330442 372068 330476 372075
rect 330229 372037 330321 372043
rect 330229 372003 330241 372037
rect 330309 372003 330321 372037
rect 330229 371997 330321 372003
rect 330505 372037 330597 372043
rect 330505 372003 330517 372037
rect 330585 372003 330597 372037
rect 330505 371997 330597 372003
rect 330626 371910 330656 372075
rect 330718 372159 330748 372172
rect 330908 372159 330942 372334
rect 330718 372147 330771 372159
rect 330718 372087 330731 372147
rect 330765 372087 330771 372147
rect 330718 372075 330771 372087
rect 330883 372147 330942 372159
rect 330883 372087 330889 372147
rect 330923 372087 330942 372147
rect 330883 372076 330942 372087
rect 330994 372159 331028 372334
rect 331057 372231 331149 372237
rect 331057 372197 331069 372231
rect 331137 372197 331149 372231
rect 331057 372191 331149 372197
rect 331333 372231 331425 372237
rect 331333 372197 331345 372231
rect 331413 372197 331425 372231
rect 331333 372191 331425 372197
rect 331180 372159 331210 372172
rect 330994 372147 331047 372159
rect 330994 372087 331007 372147
rect 331041 372087 331047 372147
rect 330883 372075 330929 372076
rect 330994 372075 331047 372087
rect 331159 372147 331210 372159
rect 331159 372087 331165 372147
rect 331199 372087 331210 372147
rect 331159 372075 331210 372087
rect 330718 371910 330748 372075
rect 330994 372072 331028 372075
rect 330781 372037 330873 372043
rect 330781 372003 330793 372037
rect 330861 372003 330873 372037
rect 330781 371997 330873 372003
rect 331057 372037 331149 372043
rect 331057 372003 331069 372037
rect 331137 372003 331149 372037
rect 331057 371997 331149 372003
rect 331180 371910 331210 372075
rect 331272 372159 331302 372172
rect 331458 372159 331492 372334
rect 331272 372147 331323 372159
rect 331272 372087 331283 372147
rect 331317 372087 331323 372147
rect 331272 372075 331323 372087
rect 331435 372147 331492 372159
rect 331435 372087 331441 372147
rect 331475 372087 331492 372147
rect 331435 372075 331492 372087
rect 331272 371910 331302 372075
rect 331458 372072 331492 372075
rect 331546 372159 331580 372334
rect 331609 372231 331701 372237
rect 331609 372197 331621 372231
rect 331689 372197 331701 372231
rect 331609 372191 331701 372197
rect 331885 372231 331977 372237
rect 331885 372197 331897 372231
rect 331965 372197 331977 372231
rect 331885 372191 331977 372197
rect 331732 372159 331762 372172
rect 331546 372147 331599 372159
rect 331546 372087 331559 372147
rect 331593 372087 331599 372147
rect 331546 372075 331599 372087
rect 331711 372147 331762 372159
rect 331711 372087 331717 372147
rect 331751 372087 331762 372147
rect 331711 372075 331762 372087
rect 331546 372070 331580 372075
rect 331333 372037 331425 372043
rect 331333 372003 331345 372037
rect 331413 372003 331425 372037
rect 331333 371997 331425 372003
rect 331609 372037 331701 372043
rect 331609 372003 331621 372037
rect 331689 372003 331701 372037
rect 331609 371997 331701 372003
rect 331732 371910 331762 372075
rect 331818 372159 331848 372172
rect 332014 372159 332048 372334
rect 331818 372147 331875 372159
rect 331818 372087 331835 372147
rect 331869 372087 331875 372147
rect 331818 372075 331875 372087
rect 331987 372147 332048 372159
rect 331987 372087 331993 372147
rect 332027 372087 332048 372147
rect 331987 372075 332048 372087
rect 331818 371910 331848 372075
rect 332014 372066 332048 372075
rect 332096 372159 332130 372334
rect 332161 372231 332253 372237
rect 332161 372197 332173 372231
rect 332241 372197 332253 372231
rect 332161 372191 332253 372197
rect 332437 372231 332529 372237
rect 332437 372197 332449 372231
rect 332517 372197 332529 372231
rect 332437 372191 332529 372197
rect 332286 372159 332316 372172
rect 332096 372147 332151 372159
rect 332096 372087 332111 372147
rect 332145 372087 332151 372147
rect 332096 372075 332151 372087
rect 332263 372147 332316 372159
rect 332263 372087 332269 372147
rect 332303 372087 332316 372147
rect 332263 372075 332316 372087
rect 332096 372072 332130 372075
rect 331885 372037 331977 372043
rect 331885 372003 331897 372037
rect 331965 372003 331977 372037
rect 331885 371997 331977 372003
rect 332161 372037 332253 372043
rect 332161 372003 332173 372037
rect 332241 372003 332253 372037
rect 332161 371997 332253 372003
rect 332286 371910 332316 372075
rect 332374 372159 332404 372170
rect 332568 372159 332602 372334
rect 332374 372147 332427 372159
rect 332374 372087 332387 372147
rect 332421 372087 332427 372147
rect 332374 372075 332427 372087
rect 332539 372147 332602 372159
rect 332539 372087 332545 372147
rect 332579 372087 332602 372147
rect 332539 372075 332602 372087
rect 332374 371910 332404 372075
rect 332568 372070 332602 372075
rect 332646 372159 332680 372334
rect 332713 372231 332805 372237
rect 332713 372197 332725 372231
rect 332793 372197 332805 372231
rect 332713 372191 332805 372197
rect 332989 372231 333081 372237
rect 332989 372197 333001 372231
rect 333069 372197 333081 372231
rect 332989 372191 333081 372197
rect 332838 372159 332868 372174
rect 332646 372147 332703 372159
rect 332646 372087 332663 372147
rect 332697 372087 332703 372147
rect 332646 372075 332703 372087
rect 332815 372147 332868 372159
rect 332815 372087 332821 372147
rect 332855 372087 332868 372147
rect 332815 372075 332868 372087
rect 332646 372072 332680 372075
rect 332437 372037 332529 372043
rect 332437 372003 332449 372037
rect 332517 372003 332529 372037
rect 332437 371997 332529 372003
rect 332713 372037 332805 372043
rect 332713 372003 332725 372037
rect 332793 372003 332805 372037
rect 332713 371997 332805 372003
rect 332838 371910 332868 372075
rect 332926 372159 332956 372174
rect 333124 372159 333158 372334
rect 332926 372147 332979 372159
rect 332926 372087 332939 372147
rect 332973 372087 332979 372147
rect 332926 372075 332979 372087
rect 333091 372147 333158 372159
rect 333091 372087 333097 372147
rect 333131 372087 333158 372147
rect 333091 372075 333158 372087
rect 332926 371910 332956 372075
rect 333124 372062 333158 372075
rect 333198 372159 333232 372334
rect 333265 372231 333357 372237
rect 333265 372197 333277 372231
rect 333345 372197 333357 372231
rect 333265 372191 333357 372197
rect 333541 372231 333633 372237
rect 333541 372197 333553 372231
rect 333621 372197 333633 372231
rect 333541 372191 333633 372197
rect 333388 372159 333418 372176
rect 333198 372147 333255 372159
rect 333198 372087 333215 372147
rect 333249 372087 333255 372147
rect 333198 372075 333255 372087
rect 333367 372147 333418 372159
rect 333367 372087 333373 372147
rect 333407 372087 333418 372147
rect 333367 372075 333418 372087
rect 333198 372066 333232 372075
rect 332989 372037 333081 372043
rect 332989 372003 333001 372037
rect 333069 372003 333081 372037
rect 332989 371997 333081 372003
rect 333265 372037 333357 372043
rect 333265 372003 333277 372037
rect 333345 372003 333357 372037
rect 333265 371997 333357 372003
rect 333388 371910 333418 372075
rect 333476 372159 333506 372174
rect 333668 372159 333702 372334
rect 333476 372147 333531 372159
rect 333476 372087 333491 372147
rect 333525 372087 333531 372147
rect 333476 372075 333531 372087
rect 333643 372147 333702 372159
rect 333643 372087 333649 372147
rect 333683 372087 333702 372147
rect 333643 372075 333702 372087
rect 333476 371910 333506 372075
rect 333668 372062 333702 372075
rect 333748 372159 333782 372334
rect 333817 372231 333909 372237
rect 333817 372197 333829 372231
rect 333897 372197 333909 372231
rect 333817 372191 333909 372197
rect 334093 372231 334185 372237
rect 334093 372197 334105 372231
rect 334173 372197 334185 372231
rect 334093 372191 334185 372197
rect 333940 372159 333970 372174
rect 333748 372147 333807 372159
rect 333748 372087 333767 372147
rect 333801 372087 333807 372147
rect 333748 372075 333807 372087
rect 333919 372147 333970 372159
rect 333919 372087 333925 372147
rect 333959 372087 333970 372147
rect 333919 372075 333970 372087
rect 333748 372060 333782 372075
rect 333541 372037 333633 372043
rect 333541 372003 333553 372037
rect 333621 372003 333633 372037
rect 333541 371997 333633 372003
rect 333817 372037 333909 372043
rect 333817 372003 333829 372037
rect 333897 372003 333909 372037
rect 333817 371997 333909 372003
rect 333940 371910 333970 372075
rect 334028 372159 334058 372176
rect 334224 372159 334258 372334
rect 334028 372147 334083 372159
rect 334028 372087 334043 372147
rect 334077 372087 334083 372147
rect 334028 372075 334083 372087
rect 334195 372147 334258 372159
rect 334195 372087 334201 372147
rect 334235 372087 334258 372147
rect 334195 372075 334258 372087
rect 334028 371910 334058 372075
rect 334224 372062 334258 372075
rect 334298 372159 334332 372334
rect 334369 372231 334461 372237
rect 334369 372197 334381 372231
rect 334449 372197 334461 372231
rect 334369 372191 334461 372197
rect 334645 372231 334737 372237
rect 334645 372197 334657 372231
rect 334725 372197 334737 372231
rect 334645 372191 334737 372197
rect 334492 372159 334522 372174
rect 334298 372147 334359 372159
rect 334298 372087 334319 372147
rect 334353 372087 334359 372147
rect 334298 372075 334359 372087
rect 334471 372147 334522 372159
rect 334471 372087 334477 372147
rect 334511 372087 334522 372147
rect 334471 372075 334522 372087
rect 334298 372060 334332 372075
rect 334093 372037 334185 372043
rect 334093 372003 334105 372037
rect 334173 372003 334185 372037
rect 334093 371997 334185 372003
rect 334369 372037 334461 372043
rect 334369 372003 334381 372037
rect 334449 372003 334461 372037
rect 334369 371997 334461 372003
rect 334492 371910 334522 372075
rect 334582 372159 334612 372176
rect 334774 372159 334808 372334
rect 334582 372147 334635 372159
rect 334582 372087 334595 372147
rect 334629 372087 334635 372147
rect 334582 372075 334635 372087
rect 334747 372147 334808 372159
rect 334747 372087 334753 372147
rect 334787 372087 334808 372147
rect 334747 372075 334808 372087
rect 334582 371910 334612 372075
rect 334774 372064 334808 372075
rect 334850 372159 334884 372334
rect 334921 372231 335013 372237
rect 334921 372197 334933 372231
rect 335001 372197 335013 372231
rect 334921 372191 335013 372197
rect 335197 372231 335289 372237
rect 335197 372197 335209 372231
rect 335277 372197 335289 372231
rect 335197 372191 335289 372197
rect 335044 372159 335074 372174
rect 334850 372147 334911 372159
rect 334850 372087 334871 372147
rect 334905 372087 334911 372147
rect 334850 372075 334911 372087
rect 335023 372147 335074 372159
rect 335023 372087 335029 372147
rect 335063 372087 335074 372147
rect 335023 372075 335074 372087
rect 334850 372064 334884 372075
rect 334645 372037 334737 372043
rect 334645 372003 334657 372037
rect 334725 372003 334737 372037
rect 334645 371997 334737 372003
rect 334921 372037 335013 372043
rect 334921 372003 334933 372037
rect 335001 372003 335013 372037
rect 334921 371997 335013 372003
rect 335044 371910 335074 372075
rect 335134 372159 335164 372176
rect 335324 372159 335358 372334
rect 335134 372147 335187 372159
rect 335134 372087 335147 372147
rect 335181 372087 335187 372147
rect 335134 372075 335187 372087
rect 335299 372147 335358 372159
rect 335299 372087 335305 372147
rect 335339 372087 335358 372147
rect 335299 372075 335358 372087
rect 335134 371910 335164 372075
rect 335324 372068 335358 372075
rect 335406 372159 335440 372334
rect 335473 372231 335565 372237
rect 335473 372197 335485 372231
rect 335553 372197 335565 372231
rect 335473 372191 335565 372197
rect 335749 372231 335841 372237
rect 335749 372197 335761 372231
rect 335829 372197 335841 372231
rect 335749 372191 335841 372197
rect 335598 372159 335628 372180
rect 335406 372147 335463 372159
rect 335406 372087 335423 372147
rect 335457 372087 335463 372147
rect 335406 372075 335463 372087
rect 335575 372147 335628 372159
rect 335575 372087 335581 372147
rect 335615 372087 335628 372147
rect 335575 372075 335628 372087
rect 335406 372066 335440 372075
rect 335197 372037 335289 372043
rect 335197 372003 335209 372037
rect 335277 372003 335289 372037
rect 335197 371997 335289 372003
rect 335473 372037 335565 372043
rect 335473 372003 335485 372037
rect 335553 372003 335565 372037
rect 335473 371997 335565 372003
rect 335598 371910 335628 372075
rect 335688 372159 335718 372182
rect 335876 372159 335910 372334
rect 335688 372147 335739 372159
rect 335688 372087 335699 372147
rect 335733 372087 335739 372147
rect 335688 372075 335739 372087
rect 335851 372147 335910 372159
rect 335851 372087 335857 372147
rect 335891 372087 335910 372147
rect 335851 372075 335910 372087
rect 335688 371910 335718 372075
rect 335876 372072 335910 372075
rect 335954 372159 335988 372334
rect 336025 372231 336117 372237
rect 336025 372197 336037 372231
rect 336105 372197 336117 372231
rect 336025 372191 336117 372197
rect 336301 372231 336393 372237
rect 336301 372197 336313 372231
rect 336381 372197 336393 372231
rect 336301 372191 336393 372197
rect 336152 372159 336182 372182
rect 335954 372147 336015 372159
rect 335954 372087 335975 372147
rect 336009 372087 336015 372147
rect 335954 372075 336015 372087
rect 336127 372147 336182 372159
rect 336127 372087 336133 372147
rect 336167 372087 336182 372147
rect 336127 372075 336182 372087
rect 335954 372074 335988 372075
rect 335749 372037 335841 372043
rect 335749 372003 335761 372037
rect 335829 372003 335841 372037
rect 335749 371997 335841 372003
rect 336025 372037 336117 372043
rect 336025 372003 336037 372037
rect 336105 372003 336117 372037
rect 336025 371997 336117 372003
rect 336152 371910 336182 372075
rect 336238 372159 336268 372186
rect 336426 372159 336460 372334
rect 336238 372147 336291 372159
rect 336238 372087 336251 372147
rect 336285 372087 336291 372147
rect 336238 372075 336291 372087
rect 336403 372147 336460 372159
rect 336403 372087 336409 372147
rect 336443 372087 336460 372147
rect 336403 372075 336460 372087
rect 336238 371910 336268 372075
rect 336426 372070 336460 372075
rect 336510 372159 336544 372334
rect 336577 372231 336669 372237
rect 336577 372197 336589 372231
rect 336657 372197 336669 372231
rect 336577 372191 336669 372197
rect 336853 372231 336945 372237
rect 336853 372197 336865 372231
rect 336933 372197 336945 372231
rect 336853 372191 336945 372197
rect 336698 372159 336728 372172
rect 336510 372147 336567 372159
rect 336510 372087 336527 372147
rect 336561 372087 336567 372147
rect 336510 372075 336567 372087
rect 336679 372147 336728 372159
rect 336679 372087 336685 372147
rect 336719 372087 336728 372147
rect 336679 372075 336728 372087
rect 336510 372068 336544 372075
rect 336301 372037 336393 372043
rect 336301 372003 336313 372037
rect 336381 372003 336393 372037
rect 336301 371997 336393 372003
rect 336577 372037 336669 372043
rect 336577 372003 336589 372037
rect 336657 372003 336669 372037
rect 336577 371997 336669 372003
rect 336698 371910 336728 372075
rect 336790 372159 336820 372170
rect 336978 372159 337012 372334
rect 336790 372147 336843 372159
rect 336790 372087 336803 372147
rect 336837 372087 336843 372147
rect 336790 372075 336843 372087
rect 336955 372147 337012 372159
rect 336955 372087 336961 372147
rect 336995 372087 337012 372147
rect 336955 372075 337012 372087
rect 336790 371910 336820 372075
rect 336978 372070 337012 372075
rect 337062 372159 337096 372334
rect 337129 372231 337221 372237
rect 337129 372197 337141 372231
rect 337209 372197 337221 372231
rect 337129 372191 337221 372197
rect 337405 372231 337497 372237
rect 337405 372197 337417 372231
rect 337485 372197 337497 372231
rect 337405 372191 337497 372197
rect 337254 372159 337284 372172
rect 337062 372147 337119 372159
rect 337062 372087 337079 372147
rect 337113 372087 337119 372147
rect 337062 372075 337119 372087
rect 337231 372147 337284 372159
rect 337231 372087 337237 372147
rect 337271 372087 337284 372147
rect 337231 372075 337284 372087
rect 337062 372072 337096 372075
rect 336853 372037 336945 372043
rect 336853 372003 336865 372037
rect 336933 372003 336945 372037
rect 336853 371997 336945 372003
rect 337129 372037 337221 372043
rect 337129 372003 337141 372037
rect 337209 372003 337221 372037
rect 337129 371997 337221 372003
rect 337254 371910 337284 372075
rect 337338 372159 337368 372172
rect 337532 372159 337566 372334
rect 337338 372147 337395 372159
rect 337338 372087 337355 372147
rect 337389 372087 337395 372147
rect 337338 372075 337395 372087
rect 337507 372147 337566 372159
rect 337507 372087 337513 372147
rect 337547 372087 337566 372147
rect 337507 372076 337566 372087
rect 337610 372159 337644 372334
rect 337681 372231 337773 372237
rect 337681 372197 337693 372231
rect 337761 372197 337773 372231
rect 337681 372191 337773 372197
rect 337804 372159 337834 372172
rect 337610 372147 337671 372159
rect 337610 372087 337631 372147
rect 337665 372087 337671 372147
rect 337507 372075 337553 372076
rect 337610 372075 337671 372087
rect 337783 372147 337834 372159
rect 337783 372087 337789 372147
rect 337823 372087 337834 372147
rect 337783 372075 337834 372087
rect 337924 372082 337958 372334
rect 337338 371910 337368 372075
rect 337610 372074 337644 372075
rect 337405 372037 337497 372043
rect 337405 372003 337417 372037
rect 337485 372003 337497 372037
rect 337405 371997 337497 372003
rect 337681 372037 337773 372043
rect 337681 372003 337693 372037
rect 337761 372003 337773 372037
rect 337681 371997 337773 372003
rect 337804 371910 337834 372075
rect 323667 371868 337836 371910
rect 337794 371866 337836 371868
rect 158318 371723 159188 371755
rect 143461 371657 159188 371723
rect 143341 371553 143433 371559
rect 143341 371519 143353 371553
rect 143421 371519 143433 371553
rect 143341 371513 143433 371519
rect 143466 371481 143506 371657
rect 143285 371469 143331 371481
rect 141258 371411 143291 371469
rect 141258 369730 142348 371411
rect 143127 371233 143169 371411
rect 143285 371409 143291 371411
rect 143325 371409 143331 371469
rect 143285 371397 143331 371409
rect 143443 371469 143506 371481
rect 143443 371409 143449 371469
rect 143483 371409 143506 371469
rect 143443 371397 143506 371409
rect 143466 371391 143506 371397
rect 143548 371481 143588 371657
rect 143617 371553 143709 371559
rect 143617 371519 143629 371553
rect 143697 371519 143709 371553
rect 143617 371513 143709 371519
rect 143893 371553 143985 371559
rect 143893 371519 143905 371553
rect 143973 371519 143985 371553
rect 143893 371513 143985 371519
rect 143742 371481 143772 371489
rect 143548 371469 143607 371481
rect 143548 371409 143567 371469
rect 143601 371409 143607 371469
rect 143548 371397 143607 371409
rect 143719 371469 143772 371481
rect 143719 371409 143725 371469
rect 143759 371409 143772 371469
rect 143719 371397 143772 371409
rect 143548 371393 143588 371397
rect 143341 371359 143433 371365
rect 143341 371325 143353 371359
rect 143421 371325 143433 371359
rect 143341 371319 143433 371325
rect 143617 371359 143709 371365
rect 143617 371325 143629 371359
rect 143697 371325 143709 371359
rect 143617 371319 143709 371325
rect 143742 371233 143772 371397
rect 143828 371481 143858 371489
rect 144024 371481 144064 371657
rect 143828 371469 143883 371481
rect 143828 371409 143843 371469
rect 143877 371409 143883 371469
rect 143828 371397 143883 371409
rect 143995 371469 144064 371481
rect 143995 371409 144001 371469
rect 144035 371409 144064 371469
rect 143995 371397 144064 371409
rect 143828 371233 143858 371397
rect 144024 371393 144064 371397
rect 144092 371481 144132 371657
rect 144169 371553 144261 371559
rect 144169 371519 144181 371553
rect 144249 371519 144261 371553
rect 144169 371513 144261 371519
rect 144445 371553 144537 371559
rect 144445 371519 144457 371553
rect 144525 371519 144537 371553
rect 144445 371513 144537 371519
rect 144296 371481 144326 371489
rect 144092 371469 144159 371481
rect 144092 371409 144119 371469
rect 144153 371409 144159 371469
rect 144092 371397 144159 371409
rect 144271 371469 144326 371481
rect 144271 371409 144277 371469
rect 144311 371409 144326 371469
rect 144271 371397 144326 371409
rect 144092 371393 144132 371397
rect 143893 371359 143985 371365
rect 143893 371325 143905 371359
rect 143973 371325 143985 371359
rect 143893 371319 143985 371325
rect 144169 371359 144261 371365
rect 144169 371325 144181 371359
rect 144249 371325 144261 371359
rect 144169 371319 144261 371325
rect 144296 371233 144326 371397
rect 144382 371481 144412 371489
rect 144572 371481 144612 371657
rect 144382 371469 144435 371481
rect 144382 371409 144395 371469
rect 144429 371409 144435 371469
rect 144382 371397 144435 371409
rect 144547 371469 144612 371481
rect 144547 371409 144553 371469
rect 144587 371409 144612 371469
rect 144547 371397 144612 371409
rect 144382 371233 144412 371397
rect 144572 371389 144612 371397
rect 144644 371481 144684 371657
rect 144721 371553 144813 371559
rect 144721 371519 144733 371553
rect 144801 371519 144813 371553
rect 144721 371513 144813 371519
rect 144997 371553 145089 371559
rect 144997 371519 145009 371553
rect 145077 371519 145089 371553
rect 144997 371513 145089 371519
rect 144844 371481 144874 371489
rect 144644 371469 144711 371481
rect 144644 371409 144671 371469
rect 144705 371409 144711 371469
rect 144644 371397 144711 371409
rect 144823 371469 144874 371481
rect 144823 371409 144829 371469
rect 144863 371409 144874 371469
rect 144823 371397 144874 371409
rect 144644 371393 144684 371397
rect 144445 371359 144537 371365
rect 144445 371325 144457 371359
rect 144525 371325 144537 371359
rect 144445 371319 144537 371325
rect 144721 371359 144813 371365
rect 144721 371325 144733 371359
rect 144801 371325 144813 371359
rect 144721 371319 144813 371325
rect 144844 371233 144874 371397
rect 144936 371481 144966 371487
rect 145124 371481 145164 371657
rect 144936 371469 144987 371481
rect 144936 371409 144947 371469
rect 144981 371409 144987 371469
rect 144936 371397 144987 371409
rect 145099 371469 145164 371481
rect 145099 371409 145105 371469
rect 145139 371409 145164 371469
rect 145099 371397 145164 371409
rect 145204 371481 145244 371657
rect 145273 371553 145365 371559
rect 145273 371519 145285 371553
rect 145353 371519 145365 371553
rect 145273 371513 145365 371519
rect 145549 371553 145641 371559
rect 145549 371519 145561 371553
rect 145629 371519 145641 371553
rect 145549 371513 145641 371519
rect 145394 371481 145424 371487
rect 145204 371469 145263 371481
rect 145204 371409 145223 371469
rect 145257 371409 145263 371469
rect 145204 371397 145263 371409
rect 145375 371469 145424 371481
rect 145375 371409 145381 371469
rect 145415 371409 145424 371469
rect 145375 371397 145424 371409
rect 144936 371233 144966 371397
rect 144997 371359 145089 371365
rect 144997 371325 145009 371359
rect 145077 371325 145089 371359
rect 144997 371319 145089 371325
rect 145273 371359 145365 371365
rect 145273 371325 145285 371359
rect 145353 371325 145365 371359
rect 145273 371319 145365 371325
rect 145394 371233 145424 371397
rect 145486 371481 145516 371485
rect 145678 371481 145718 371657
rect 145486 371469 145539 371481
rect 145486 371409 145499 371469
rect 145533 371409 145539 371469
rect 145486 371397 145539 371409
rect 145651 371469 145718 371481
rect 145651 371409 145657 371469
rect 145691 371409 145718 371469
rect 145651 371397 145718 371409
rect 145486 371233 145516 371397
rect 145678 371393 145718 371397
rect 145752 371481 145792 371657
rect 145825 371553 145917 371559
rect 145825 371519 145837 371553
rect 145905 371519 145917 371553
rect 145825 371513 145917 371519
rect 146101 371553 146193 371559
rect 146101 371519 146113 371553
rect 146181 371519 146193 371553
rect 146101 371513 146193 371519
rect 145950 371481 145980 371485
rect 145752 371469 145815 371481
rect 145752 371409 145775 371469
rect 145809 371409 145815 371469
rect 145752 371397 145815 371409
rect 145927 371469 145980 371481
rect 145927 371409 145933 371469
rect 145967 371409 145980 371469
rect 145927 371397 145980 371409
rect 145752 371395 145792 371397
rect 145549 371359 145641 371365
rect 145549 371325 145561 371359
rect 145629 371325 145641 371359
rect 145549 371319 145641 371325
rect 145825 371359 145917 371365
rect 145825 371325 145837 371359
rect 145905 371325 145917 371359
rect 145825 371319 145917 371325
rect 145950 371233 145980 371397
rect 146038 371481 146068 371483
rect 146230 371481 146270 371657
rect 146038 371469 146091 371481
rect 146038 371409 146051 371469
rect 146085 371409 146091 371469
rect 146038 371397 146091 371409
rect 146203 371469 146270 371481
rect 146203 371409 146209 371469
rect 146243 371409 146270 371469
rect 146203 371397 146270 371409
rect 146038 371233 146068 371397
rect 146230 371391 146270 371397
rect 146300 371481 146340 371657
rect 146377 371553 146469 371559
rect 146377 371519 146389 371553
rect 146457 371519 146469 371553
rect 146377 371513 146469 371519
rect 146653 371553 146745 371559
rect 146653 371519 146665 371553
rect 146733 371519 146745 371553
rect 146653 371513 146745 371519
rect 146500 371481 146530 371483
rect 146300 371469 146367 371481
rect 146300 371409 146327 371469
rect 146361 371409 146367 371469
rect 146300 371397 146367 371409
rect 146479 371469 146530 371481
rect 146479 371409 146485 371469
rect 146519 371409 146530 371469
rect 146479 371397 146530 371409
rect 146300 371395 146340 371397
rect 146101 371359 146193 371365
rect 146377 371363 146469 371365
rect 146101 371325 146113 371359
rect 146181 371325 146193 371359
rect 146374 371359 146469 371363
rect 146374 371330 146389 371359
rect 146101 371319 146193 371325
rect 146377 371325 146389 371330
rect 146457 371325 146469 371359
rect 146377 371319 146469 371325
rect 146500 371233 146530 371397
rect 146588 371481 146618 371483
rect 146778 371481 146818 371657
rect 146588 371469 146643 371481
rect 146588 371409 146603 371469
rect 146637 371409 146643 371469
rect 146588 371397 146643 371409
rect 146755 371469 146818 371481
rect 146755 371409 146761 371469
rect 146795 371409 146818 371469
rect 146755 371397 146818 371409
rect 146588 371233 146618 371397
rect 146778 371391 146818 371397
rect 146856 371481 146896 371657
rect 146929 371553 147021 371559
rect 146929 371519 146941 371553
rect 147009 371519 147021 371553
rect 146929 371513 147021 371519
rect 147205 371553 147297 371559
rect 147205 371519 147217 371553
rect 147285 371519 147297 371553
rect 147205 371513 147297 371519
rect 147052 371481 147082 371485
rect 146856 371469 146919 371481
rect 146856 371409 146879 371469
rect 146913 371409 146919 371469
rect 146856 371397 146919 371409
rect 147031 371469 147082 371481
rect 147031 371409 147037 371469
rect 147071 371409 147082 371469
rect 147031 371397 147082 371409
rect 146856 371395 146896 371397
rect 146653 371359 146745 371365
rect 146653 371325 146665 371359
rect 146733 371325 146745 371359
rect 146653 371319 146745 371325
rect 146929 371359 147021 371365
rect 146929 371325 146941 371359
rect 147009 371325 147021 371359
rect 146929 371319 147021 371325
rect 147052 371233 147082 371397
rect 147140 371481 147170 371485
rect 147332 371481 147372 371657
rect 147140 371469 147195 371481
rect 147140 371409 147155 371469
rect 147189 371409 147195 371469
rect 147140 371397 147195 371409
rect 147307 371469 147372 371481
rect 147307 371409 147313 371469
rect 147347 371409 147372 371469
rect 147307 371397 147372 371409
rect 147140 371233 147170 371397
rect 147332 371383 147372 371397
rect 147410 371481 147450 371657
rect 147481 371553 147573 371559
rect 147481 371519 147493 371553
rect 147561 371519 147573 371553
rect 147481 371513 147573 371519
rect 147757 371553 147849 371559
rect 147757 371519 147769 371553
rect 147837 371519 147849 371553
rect 147757 371513 147849 371519
rect 147604 371481 147634 371485
rect 147410 371469 147471 371481
rect 147410 371409 147431 371469
rect 147465 371409 147471 371469
rect 147410 371397 147471 371409
rect 147583 371469 147634 371481
rect 147583 371409 147589 371469
rect 147623 371409 147634 371469
rect 147583 371397 147634 371409
rect 147410 371391 147450 371397
rect 147205 371359 147297 371365
rect 147205 371325 147217 371359
rect 147285 371325 147297 371359
rect 147205 371319 147297 371325
rect 147481 371359 147573 371365
rect 147481 371325 147493 371359
rect 147561 371325 147573 371359
rect 147481 371319 147573 371325
rect 147604 371233 147634 371397
rect 147696 371481 147726 371485
rect 147888 371481 147928 371657
rect 147696 371469 147747 371481
rect 147696 371409 147707 371469
rect 147741 371409 147747 371469
rect 147696 371397 147747 371409
rect 147859 371469 147928 371481
rect 147859 371409 147865 371469
rect 147899 371409 147928 371469
rect 147859 371397 147928 371409
rect 147962 371481 148002 371657
rect 148033 371553 148125 371559
rect 148033 371519 148045 371553
rect 148113 371519 148125 371553
rect 148033 371513 148125 371519
rect 148309 371553 148401 371559
rect 148309 371519 148321 371553
rect 148389 371519 148401 371553
rect 148309 371513 148401 371519
rect 148158 371481 148188 371495
rect 147962 371469 148023 371481
rect 147962 371409 147983 371469
rect 148017 371409 148023 371469
rect 147962 371397 148023 371409
rect 148135 371469 148188 371481
rect 148135 371409 148141 371469
rect 148175 371409 148188 371469
rect 148135 371397 148188 371409
rect 147696 371233 147726 371397
rect 147888 371393 147928 371397
rect 147757 371359 147849 371365
rect 147757 371325 147769 371359
rect 147837 371325 147849 371359
rect 147757 371319 147849 371325
rect 148033 371359 148125 371365
rect 148033 371325 148045 371359
rect 148113 371325 148125 371359
rect 148033 371319 148125 371325
rect 148158 371233 148188 371397
rect 148244 371481 148274 371493
rect 148432 371481 148466 371657
rect 148244 371469 148299 371481
rect 148244 371409 148259 371469
rect 148293 371409 148299 371469
rect 148244 371397 148299 371409
rect 148411 371469 148466 371481
rect 148411 371409 148417 371469
rect 148451 371409 148466 371469
rect 148411 371397 148466 371409
rect 148244 371233 148274 371397
rect 148432 371393 148466 371397
rect 148522 371481 148556 371657
rect 148585 371553 148677 371559
rect 148585 371519 148597 371553
rect 148665 371519 148677 371553
rect 148585 371513 148677 371519
rect 148861 371553 148953 371559
rect 148861 371519 148873 371553
rect 148941 371519 148953 371553
rect 148861 371513 148953 371519
rect 148712 371481 148742 371491
rect 148522 371469 148575 371481
rect 148522 371409 148535 371469
rect 148569 371409 148575 371469
rect 148522 371397 148575 371409
rect 148687 371469 148742 371481
rect 148687 371409 148693 371469
rect 148727 371409 148742 371469
rect 148687 371397 148742 371409
rect 148522 371393 148556 371397
rect 148309 371359 148401 371365
rect 148309 371325 148321 371359
rect 148389 371325 148401 371359
rect 148309 371319 148401 371325
rect 148585 371359 148677 371365
rect 148585 371325 148597 371359
rect 148665 371325 148677 371359
rect 148585 371319 148677 371325
rect 148712 371233 148742 371397
rect 148798 371481 148828 371491
rect 148988 371481 149022 371657
rect 148798 371469 148851 371481
rect 148798 371409 148811 371469
rect 148845 371409 148851 371469
rect 148798 371397 148851 371409
rect 148963 371469 149022 371481
rect 148963 371409 148969 371469
rect 149003 371409 149022 371469
rect 148963 371397 149022 371409
rect 149072 371481 149106 371657
rect 149137 371553 149229 371559
rect 149137 371519 149149 371553
rect 149217 371519 149229 371553
rect 149137 371513 149229 371519
rect 149264 371481 149298 371495
rect 149072 371469 149127 371481
rect 149072 371409 149087 371469
rect 149121 371409 149127 371469
rect 149072 371397 149127 371409
rect 149239 371469 149298 371481
rect 149239 371409 149245 371469
rect 149279 371409 149298 371469
rect 149239 371397 149298 371409
rect 148798 371233 148828 371397
rect 148988 371393 149022 371397
rect 148861 371359 148953 371365
rect 148861 371325 148873 371359
rect 148941 371325 148953 371359
rect 148861 371319 148953 371325
rect 149137 371359 149229 371365
rect 149137 371325 149149 371359
rect 149217 371325 149229 371359
rect 149137 371319 149229 371325
rect 149264 371233 149298 371397
rect 149346 371481 149380 371657
rect 149413 371553 149505 371559
rect 149413 371519 149425 371553
rect 149493 371519 149505 371553
rect 149413 371513 149505 371519
rect 149689 371553 149781 371559
rect 149689 371519 149701 371553
rect 149769 371519 149781 371553
rect 149689 371513 149781 371519
rect 149538 371481 149568 371493
rect 149346 371469 149403 371481
rect 149346 371409 149363 371469
rect 149397 371409 149403 371469
rect 149346 371397 149403 371409
rect 149515 371469 149568 371481
rect 149515 371409 149521 371469
rect 149555 371409 149568 371469
rect 149515 371397 149568 371409
rect 149346 371395 149380 371397
rect 149413 371359 149505 371365
rect 149413 371325 149425 371359
rect 149493 371325 149505 371359
rect 149413 371319 149505 371325
rect 149538 371233 149568 371397
rect 149626 371481 149656 371495
rect 149816 371481 149850 371657
rect 149626 371469 149679 371481
rect 149626 371409 149639 371469
rect 149673 371409 149679 371469
rect 149626 371397 149679 371409
rect 149791 371469 149850 371481
rect 149791 371409 149797 371469
rect 149831 371409 149850 371469
rect 149791 371397 149850 371409
rect 149902 371481 149936 371657
rect 149974 371595 150189 371605
rect 149974 371559 150104 371595
rect 149965 371553 150104 371559
rect 149965 371519 149977 371553
rect 150045 371535 150104 371553
rect 150164 371535 150189 371595
rect 150045 371525 150189 371535
rect 150241 371553 150333 371559
rect 150045 371519 150057 371525
rect 149965 371513 150057 371519
rect 150241 371519 150253 371553
rect 150321 371519 150333 371553
rect 150241 371513 150333 371519
rect 150086 371481 150116 371495
rect 149902 371469 149955 371481
rect 149902 371409 149915 371469
rect 149949 371409 149955 371469
rect 149902 371397 149955 371409
rect 150067 371469 150116 371481
rect 150067 371409 150073 371469
rect 150107 371409 150116 371469
rect 150067 371397 150116 371409
rect 149626 371233 149656 371397
rect 149902 371391 149936 371397
rect 149689 371359 149781 371365
rect 149689 371325 149701 371359
rect 149769 371325 149781 371359
rect 149965 371359 150057 371365
rect 149965 371340 149977 371359
rect 149689 371319 149781 371325
rect 149829 371335 149977 371340
rect 149829 371280 149839 371335
rect 149904 371325 149977 371335
rect 150045 371325 150057 371359
rect 149904 371319 150057 371325
rect 149904 371290 150044 371319
rect 149904 371280 149914 371290
rect 149829 371275 149914 371280
rect 150086 371233 150116 371397
rect 150178 371481 150208 371495
rect 150368 371481 150402 371657
rect 150178 371469 150231 371481
rect 150178 371409 150191 371469
rect 150225 371409 150231 371469
rect 150178 371397 150231 371409
rect 150343 371469 150402 371481
rect 150343 371409 150349 371469
rect 150383 371409 150402 371469
rect 150343 371399 150402 371409
rect 150454 371481 150488 371657
rect 150517 371553 150609 371559
rect 150517 371519 150529 371553
rect 150597 371519 150609 371553
rect 150517 371513 150609 371519
rect 150793 371553 150885 371559
rect 150793 371519 150805 371553
rect 150873 371519 150885 371553
rect 150793 371513 150885 371519
rect 150640 371481 150670 371495
rect 150454 371469 150507 371481
rect 150454 371409 150467 371469
rect 150501 371409 150507 371469
rect 150343 371397 150389 371399
rect 150454 371397 150507 371409
rect 150619 371469 150670 371481
rect 150619 371409 150625 371469
rect 150659 371409 150670 371469
rect 150619 371397 150670 371409
rect 150178 371233 150208 371397
rect 150454 371395 150488 371397
rect 150241 371359 150333 371365
rect 150241 371325 150253 371359
rect 150321 371325 150333 371359
rect 150241 371319 150333 371325
rect 150517 371359 150609 371365
rect 150517 371325 150529 371359
rect 150597 371325 150609 371359
rect 150517 371319 150609 371325
rect 150640 371233 150670 371397
rect 150732 371481 150762 371495
rect 150918 371481 150952 371657
rect 150732 371469 150783 371481
rect 150732 371409 150743 371469
rect 150777 371409 150783 371469
rect 150732 371397 150783 371409
rect 150895 371469 150952 371481
rect 150895 371409 150901 371469
rect 150935 371409 150952 371469
rect 150895 371397 150952 371409
rect 150732 371233 150762 371397
rect 150918 371395 150952 371397
rect 151006 371481 151040 371657
rect 151069 371553 151161 371559
rect 151069 371519 151081 371553
rect 151149 371519 151161 371553
rect 151069 371513 151161 371519
rect 151345 371553 151437 371559
rect 151345 371519 151357 371553
rect 151425 371519 151437 371553
rect 151345 371513 151437 371519
rect 151192 371481 151222 371495
rect 151006 371469 151059 371481
rect 151006 371409 151019 371469
rect 151053 371409 151059 371469
rect 151006 371397 151059 371409
rect 151171 371469 151222 371481
rect 151171 371409 151177 371469
rect 151211 371409 151222 371469
rect 151171 371397 151222 371409
rect 151006 371393 151040 371397
rect 150793 371359 150885 371365
rect 150793 371325 150805 371359
rect 150873 371325 150885 371359
rect 150793 371319 150885 371325
rect 151069 371359 151161 371365
rect 151069 371325 151081 371359
rect 151149 371325 151161 371359
rect 151069 371319 151161 371325
rect 151192 371233 151222 371397
rect 151278 371481 151308 371495
rect 151474 371481 151508 371657
rect 151278 371469 151335 371481
rect 151278 371409 151295 371469
rect 151329 371409 151335 371469
rect 151278 371397 151335 371409
rect 151447 371469 151508 371481
rect 151447 371409 151453 371469
rect 151487 371409 151508 371469
rect 151447 371397 151508 371409
rect 151278 371233 151308 371397
rect 151474 371389 151508 371397
rect 151556 371481 151590 371657
rect 151621 371553 151713 371559
rect 151621 371519 151633 371553
rect 151701 371519 151713 371553
rect 151621 371513 151713 371519
rect 151897 371553 151989 371559
rect 151897 371519 151909 371553
rect 151977 371519 151989 371553
rect 151897 371513 151989 371519
rect 151746 371481 151776 371495
rect 151556 371469 151611 371481
rect 151556 371409 151571 371469
rect 151605 371409 151611 371469
rect 151556 371397 151611 371409
rect 151723 371469 151776 371481
rect 151723 371409 151729 371469
rect 151763 371409 151776 371469
rect 151723 371397 151776 371409
rect 151556 371395 151590 371397
rect 151345 371359 151437 371365
rect 151345 371325 151357 371359
rect 151425 371325 151437 371359
rect 151345 371319 151437 371325
rect 151621 371359 151713 371365
rect 151621 371325 151633 371359
rect 151701 371325 151713 371359
rect 151621 371319 151713 371325
rect 151746 371233 151776 371397
rect 151834 371481 151864 371493
rect 152028 371481 152062 371657
rect 151834 371469 151887 371481
rect 151834 371409 151847 371469
rect 151881 371409 151887 371469
rect 151834 371397 151887 371409
rect 151999 371469 152062 371481
rect 151999 371409 152005 371469
rect 152039 371409 152062 371469
rect 151999 371397 152062 371409
rect 151834 371233 151864 371397
rect 152028 371393 152062 371397
rect 152106 371481 152140 371657
rect 152173 371553 152265 371559
rect 152173 371519 152185 371553
rect 152253 371519 152265 371553
rect 152173 371513 152265 371519
rect 152449 371553 152541 371559
rect 152449 371519 152461 371553
rect 152529 371519 152541 371553
rect 152449 371513 152541 371519
rect 152298 371481 152328 371497
rect 152106 371469 152163 371481
rect 152106 371409 152123 371469
rect 152157 371409 152163 371469
rect 152106 371397 152163 371409
rect 152275 371469 152328 371481
rect 152275 371409 152281 371469
rect 152315 371409 152328 371469
rect 152275 371397 152328 371409
rect 152106 371395 152140 371397
rect 151897 371359 151989 371365
rect 151897 371325 151909 371359
rect 151977 371325 151989 371359
rect 151897 371319 151989 371325
rect 152173 371359 152265 371365
rect 152173 371325 152185 371359
rect 152253 371325 152265 371359
rect 152173 371319 152265 371325
rect 152298 371233 152328 371397
rect 152386 371481 152416 371497
rect 152584 371481 152618 371657
rect 152386 371469 152439 371481
rect 152386 371409 152399 371469
rect 152433 371409 152439 371469
rect 152386 371397 152439 371409
rect 152551 371469 152618 371481
rect 152551 371409 152557 371469
rect 152591 371409 152618 371469
rect 152551 371397 152618 371409
rect 152386 371233 152416 371397
rect 152584 371385 152618 371397
rect 152658 371481 152692 371657
rect 152725 371553 152817 371559
rect 152725 371519 152737 371553
rect 152805 371519 152817 371553
rect 152725 371513 152817 371519
rect 153001 371553 153093 371559
rect 153001 371519 153013 371553
rect 153081 371519 153093 371553
rect 153001 371513 153093 371519
rect 152848 371481 152878 371499
rect 152658 371469 152715 371481
rect 152658 371409 152675 371469
rect 152709 371409 152715 371469
rect 152658 371397 152715 371409
rect 152827 371469 152878 371481
rect 152827 371409 152833 371469
rect 152867 371409 152878 371469
rect 152827 371397 152878 371409
rect 152658 371389 152692 371397
rect 152449 371359 152541 371365
rect 152449 371325 152461 371359
rect 152529 371325 152541 371359
rect 152449 371319 152541 371325
rect 152725 371359 152817 371365
rect 152725 371325 152737 371359
rect 152805 371325 152817 371359
rect 152725 371319 152817 371325
rect 152848 371233 152878 371397
rect 152936 371481 152966 371497
rect 153128 371481 153162 371657
rect 152936 371469 152991 371481
rect 152936 371409 152951 371469
rect 152985 371409 152991 371469
rect 152936 371397 152991 371409
rect 153103 371469 153162 371481
rect 153103 371409 153109 371469
rect 153143 371409 153162 371469
rect 153103 371397 153162 371409
rect 152936 371233 152966 371397
rect 153128 371385 153162 371397
rect 153208 371481 153242 371657
rect 153277 371553 153369 371559
rect 153277 371519 153289 371553
rect 153357 371519 153369 371553
rect 153277 371513 153369 371519
rect 153553 371553 153645 371559
rect 153553 371519 153565 371553
rect 153633 371519 153645 371553
rect 153553 371513 153645 371519
rect 153400 371481 153430 371497
rect 153208 371469 153267 371481
rect 153208 371409 153227 371469
rect 153261 371409 153267 371469
rect 153208 371397 153267 371409
rect 153379 371469 153430 371481
rect 153379 371409 153385 371469
rect 153419 371409 153430 371469
rect 153379 371397 153430 371409
rect 153208 371383 153242 371397
rect 153001 371359 153093 371365
rect 153001 371325 153013 371359
rect 153081 371325 153093 371359
rect 153001 371319 153093 371325
rect 153277 371359 153369 371365
rect 153277 371325 153289 371359
rect 153357 371325 153369 371359
rect 153277 371319 153369 371325
rect 153400 371233 153430 371397
rect 153488 371481 153518 371499
rect 153684 371481 153718 371657
rect 153488 371469 153543 371481
rect 153488 371409 153503 371469
rect 153537 371409 153543 371469
rect 153488 371397 153543 371409
rect 153655 371469 153718 371481
rect 153655 371409 153661 371469
rect 153695 371409 153718 371469
rect 153655 371397 153718 371409
rect 153488 371233 153518 371397
rect 153684 371385 153718 371397
rect 153758 371481 153792 371657
rect 153829 371553 153921 371559
rect 153829 371519 153841 371553
rect 153909 371519 153921 371553
rect 153829 371513 153921 371519
rect 154105 371553 154197 371559
rect 154105 371519 154117 371553
rect 154185 371519 154197 371553
rect 154105 371513 154197 371519
rect 153952 371481 153982 371497
rect 153758 371469 153819 371481
rect 153758 371409 153779 371469
rect 153813 371409 153819 371469
rect 153758 371397 153819 371409
rect 153931 371469 153982 371481
rect 153931 371409 153937 371469
rect 153971 371409 153982 371469
rect 153931 371397 153982 371409
rect 153758 371383 153792 371397
rect 153553 371359 153645 371365
rect 153553 371325 153565 371359
rect 153633 371325 153645 371359
rect 153553 371319 153645 371325
rect 153829 371359 153921 371365
rect 153829 371325 153841 371359
rect 153909 371325 153921 371359
rect 153829 371319 153921 371325
rect 153952 371233 153982 371397
rect 154042 371481 154072 371499
rect 154234 371481 154268 371657
rect 154042 371469 154095 371481
rect 154042 371409 154055 371469
rect 154089 371409 154095 371469
rect 154042 371397 154095 371409
rect 154207 371469 154268 371481
rect 154207 371409 154213 371469
rect 154247 371409 154268 371469
rect 154207 371397 154268 371409
rect 154042 371233 154072 371397
rect 154234 371387 154268 371397
rect 154310 371481 154344 371657
rect 154381 371553 154473 371559
rect 154381 371519 154393 371553
rect 154461 371519 154473 371553
rect 154381 371513 154473 371519
rect 154657 371553 154749 371559
rect 154657 371519 154669 371553
rect 154737 371519 154749 371553
rect 154657 371513 154749 371519
rect 154504 371481 154534 371497
rect 154310 371469 154371 371481
rect 154310 371409 154331 371469
rect 154365 371409 154371 371469
rect 154310 371397 154371 371409
rect 154483 371469 154534 371481
rect 154483 371409 154489 371469
rect 154523 371409 154534 371469
rect 154483 371397 154534 371409
rect 154310 371387 154344 371397
rect 154105 371359 154197 371365
rect 154105 371325 154117 371359
rect 154185 371325 154197 371359
rect 154105 371319 154197 371325
rect 154381 371359 154473 371365
rect 154381 371325 154393 371359
rect 154461 371325 154473 371359
rect 154381 371319 154473 371325
rect 154504 371233 154534 371397
rect 154594 371481 154624 371499
rect 154784 371481 154818 371657
rect 154594 371469 154647 371481
rect 154594 371409 154607 371469
rect 154641 371409 154647 371469
rect 154594 371397 154647 371409
rect 154759 371469 154818 371481
rect 154759 371409 154765 371469
rect 154799 371409 154818 371469
rect 154759 371397 154818 371409
rect 154594 371233 154624 371397
rect 154784 371391 154818 371397
rect 154866 371481 154900 371657
rect 154933 371553 155025 371559
rect 154933 371519 154945 371553
rect 155013 371519 155025 371553
rect 154933 371513 155025 371519
rect 155209 371553 155301 371559
rect 155209 371519 155221 371553
rect 155289 371519 155301 371553
rect 155209 371513 155301 371519
rect 155058 371481 155088 371503
rect 154866 371469 154923 371481
rect 154866 371409 154883 371469
rect 154917 371409 154923 371469
rect 154866 371397 154923 371409
rect 155035 371469 155088 371481
rect 155035 371409 155041 371469
rect 155075 371409 155088 371469
rect 155035 371397 155088 371409
rect 154866 371389 154900 371397
rect 154657 371359 154749 371365
rect 154657 371325 154669 371359
rect 154737 371325 154749 371359
rect 154657 371319 154749 371325
rect 154933 371359 155025 371365
rect 154933 371325 154945 371359
rect 155013 371325 155025 371359
rect 154933 371319 155025 371325
rect 155058 371233 155088 371397
rect 155148 371481 155178 371505
rect 155336 371481 155370 371657
rect 155148 371469 155199 371481
rect 155148 371409 155159 371469
rect 155193 371409 155199 371469
rect 155148 371397 155199 371409
rect 155311 371469 155370 371481
rect 155311 371409 155317 371469
rect 155351 371409 155370 371469
rect 155311 371397 155370 371409
rect 155414 371481 155448 371657
rect 155485 371553 155577 371559
rect 155485 371519 155497 371553
rect 155565 371519 155577 371553
rect 155485 371513 155577 371519
rect 155761 371553 155853 371559
rect 155761 371519 155773 371553
rect 155841 371519 155853 371553
rect 155761 371513 155853 371519
rect 155612 371481 155642 371505
rect 155414 371469 155475 371481
rect 155414 371409 155435 371469
rect 155469 371409 155475 371469
rect 155414 371397 155475 371409
rect 155587 371469 155642 371481
rect 155587 371409 155593 371469
rect 155627 371409 155642 371469
rect 155587 371397 155642 371409
rect 155148 371233 155178 371397
rect 155336 371395 155370 371397
rect 155209 371359 155301 371365
rect 155209 371325 155221 371359
rect 155289 371325 155301 371359
rect 155209 371319 155301 371325
rect 155485 371359 155577 371365
rect 155485 371325 155497 371359
rect 155565 371325 155577 371359
rect 155485 371319 155577 371325
rect 155612 371233 155642 371397
rect 155698 371481 155728 371509
rect 155886 371481 155920 371657
rect 155698 371469 155751 371481
rect 155698 371409 155711 371469
rect 155745 371409 155751 371469
rect 155698 371397 155751 371409
rect 155863 371469 155920 371481
rect 155863 371409 155869 371469
rect 155903 371409 155920 371469
rect 155863 371397 155920 371409
rect 155698 371233 155728 371397
rect 155886 371393 155920 371397
rect 155970 371481 156004 371657
rect 156037 371553 156129 371559
rect 156037 371519 156049 371553
rect 156117 371519 156129 371553
rect 156037 371513 156129 371519
rect 156313 371553 156405 371559
rect 156313 371519 156325 371553
rect 156393 371519 156405 371553
rect 156313 371513 156405 371519
rect 156158 371481 156188 371495
rect 155970 371469 156027 371481
rect 155970 371409 155987 371469
rect 156021 371409 156027 371469
rect 155970 371397 156027 371409
rect 156139 371469 156188 371481
rect 156139 371409 156145 371469
rect 156179 371409 156188 371469
rect 156139 371397 156188 371409
rect 155970 371391 156004 371397
rect 155761 371359 155853 371365
rect 155761 371325 155773 371359
rect 155841 371325 155853 371359
rect 155761 371319 155853 371325
rect 156037 371359 156129 371365
rect 156037 371325 156049 371359
rect 156117 371325 156129 371359
rect 156037 371319 156129 371325
rect 156158 371233 156188 371397
rect 156250 371481 156280 371493
rect 156438 371481 156472 371657
rect 156250 371469 156303 371481
rect 156250 371409 156263 371469
rect 156297 371409 156303 371469
rect 156250 371397 156303 371409
rect 156415 371469 156472 371481
rect 156415 371409 156421 371469
rect 156455 371409 156472 371469
rect 156415 371397 156472 371409
rect 156250 371233 156280 371397
rect 156438 371393 156472 371397
rect 156522 371481 156556 371657
rect 156589 371553 156681 371559
rect 156589 371519 156601 371553
rect 156669 371519 156681 371553
rect 156589 371513 156681 371519
rect 156865 371553 156957 371559
rect 156865 371519 156877 371553
rect 156945 371519 156957 371553
rect 156865 371513 156957 371519
rect 156714 371481 156744 371495
rect 156522 371469 156579 371481
rect 156522 371409 156539 371469
rect 156573 371409 156579 371469
rect 156522 371397 156579 371409
rect 156691 371469 156744 371481
rect 156691 371409 156697 371469
rect 156731 371409 156744 371469
rect 156691 371397 156744 371409
rect 156522 371395 156556 371397
rect 156313 371359 156405 371365
rect 156313 371325 156325 371359
rect 156393 371325 156405 371359
rect 156313 371319 156405 371325
rect 156589 371359 156681 371365
rect 156589 371325 156601 371359
rect 156669 371325 156681 371359
rect 156589 371319 156681 371325
rect 156714 371233 156744 371397
rect 156798 371481 156828 371495
rect 156992 371481 157026 371657
rect 156798 371469 156855 371481
rect 156798 371409 156815 371469
rect 156849 371409 156855 371469
rect 156798 371397 156855 371409
rect 156967 371469 157026 371481
rect 156967 371409 156973 371469
rect 157007 371409 157026 371469
rect 156967 371399 157026 371409
rect 157070 371481 157104 371657
rect 157141 371553 157233 371559
rect 157141 371519 157153 371553
rect 157221 371519 157233 371553
rect 157141 371513 157233 371519
rect 157264 371481 157294 371495
rect 157070 371469 157131 371481
rect 157070 371409 157091 371469
rect 157125 371409 157131 371469
rect 156967 371397 157013 371399
rect 157070 371397 157131 371409
rect 157243 371469 157294 371481
rect 157243 371409 157249 371469
rect 157283 371409 157294 371469
rect 157243 371397 157294 371409
rect 157384 371405 157418 371657
rect 156798 371233 156828 371397
rect 156865 371359 156957 371365
rect 156865 371325 156877 371359
rect 156945 371325 156957 371359
rect 156865 371319 156957 371325
rect 157141 371359 157233 371365
rect 157141 371325 157153 371359
rect 157221 371325 157233 371359
rect 157141 371319 157233 371325
rect 157264 371233 157294 371397
rect 143127 371191 157296 371233
rect 157254 371189 157296 371191
rect 147306 371085 147446 371097
rect 147306 371029 147346 371085
rect 147424 371029 147446 371085
rect 147306 370415 147446 371029
rect 158318 370600 159188 371657
rect 230433 370873 231381 371842
rect 327846 371762 327986 371774
rect 323888 371686 323972 371718
rect 323888 371644 323904 371686
rect 323958 371644 323972 371686
rect 323888 371556 323972 371644
rect 323888 371500 323896 371556
rect 323964 371500 323972 371556
rect 323888 371492 323972 371500
rect 327846 371706 327886 371762
rect 327964 371706 327986 371762
rect 247608 371127 249092 371157
rect 232818 371061 249092 371127
rect 327846 371092 327986 371706
rect 338790 371610 339590 372334
rect 420002 372392 420088 372592
rect 420002 372328 420008 372392
rect 420080 372328 420088 372392
rect 420002 372302 420088 372328
rect 508478 372100 508924 372104
rect 508118 372060 508924 372100
rect 419006 371996 422804 372050
rect 418891 371843 418983 371849
rect 417964 371786 418164 371834
rect 418891 371809 418903 371843
rect 418971 371809 418983 371843
rect 418891 371803 418983 371809
rect 417964 371684 417996 371786
rect 418146 371684 418164 371786
rect 417964 371634 418164 371684
rect 418828 371771 418860 371788
rect 419012 371771 419042 371996
rect 418828 371759 418881 371771
rect 418828 371699 418841 371759
rect 418875 371699 418881 371759
rect 418828 371687 418881 371699
rect 418993 371759 419042 371771
rect 418993 371699 418999 371759
rect 419033 371699 419042 371759
rect 418993 371687 419042 371699
rect 338790 371364 338860 371610
rect 339000 371364 339590 371610
rect 418039 371434 418085 371634
rect 418828 371434 418860 371687
rect 419012 371666 419042 371687
rect 419102 371771 419132 371996
rect 419167 371843 419259 371849
rect 419167 371809 419179 371843
rect 419247 371809 419259 371843
rect 419167 371803 419259 371809
rect 419443 371843 419535 371849
rect 419443 371809 419455 371843
rect 419523 371809 419535 371843
rect 419443 371803 419535 371809
rect 419294 371771 419326 371790
rect 419102 371759 419157 371771
rect 419102 371699 419117 371759
rect 419151 371699 419157 371759
rect 419102 371687 419157 371699
rect 419269 371759 419326 371771
rect 419269 371699 419275 371759
rect 419309 371699 419326 371759
rect 419269 371687 419326 371699
rect 419102 371666 419132 371687
rect 418891 371649 418983 371655
rect 418891 371615 418903 371649
rect 418971 371615 418983 371649
rect 418891 371609 418983 371615
rect 419167 371649 419259 371655
rect 419167 371615 419179 371649
rect 419247 371615 419259 371649
rect 419167 371609 419259 371615
rect 419294 371434 419326 371687
rect 419376 371771 419408 371790
rect 419564 371771 419594 371996
rect 419376 371759 419433 371771
rect 419376 371699 419393 371759
rect 419427 371699 419433 371759
rect 419376 371687 419433 371699
rect 419545 371759 419594 371771
rect 419545 371699 419551 371759
rect 419585 371699 419594 371759
rect 419545 371687 419594 371699
rect 419376 371434 419408 371687
rect 419564 371668 419594 371687
rect 419654 371771 419684 371996
rect 420006 371872 420086 371882
rect 420006 371849 420008 371872
rect 419719 371843 419811 371849
rect 419719 371809 419731 371843
rect 419799 371809 419811 371843
rect 419719 371803 419811 371809
rect 419995 371843 420008 371849
rect 420076 371849 420086 371872
rect 419995 371809 420007 371843
rect 420076 371816 420087 371849
rect 420075 371809 420087 371816
rect 419995 371803 420087 371809
rect 419846 371771 419878 371790
rect 419654 371759 419709 371771
rect 419654 371699 419669 371759
rect 419703 371699 419709 371759
rect 419654 371687 419709 371699
rect 419821 371759 419878 371771
rect 419821 371699 419827 371759
rect 419861 371699 419878 371759
rect 419821 371687 419878 371699
rect 419654 371666 419684 371687
rect 419443 371649 419535 371655
rect 419443 371615 419455 371649
rect 419523 371615 419535 371649
rect 419443 371609 419535 371615
rect 419719 371649 419811 371655
rect 419719 371615 419731 371649
rect 419799 371615 419811 371649
rect 419719 371609 419811 371615
rect 419846 371434 419878 371687
rect 419934 371771 419966 371788
rect 420118 371771 420148 371996
rect 419934 371759 419985 371771
rect 419934 371699 419945 371759
rect 419979 371699 419985 371759
rect 419934 371687 419985 371699
rect 420097 371759 420148 371771
rect 420097 371699 420103 371759
rect 420137 371699 420148 371759
rect 420097 371687 420148 371699
rect 419934 371434 419966 371687
rect 420118 371662 420148 371687
rect 420208 371771 420238 371996
rect 420271 371843 420363 371849
rect 420271 371809 420283 371843
rect 420351 371809 420363 371843
rect 420271 371803 420363 371809
rect 420547 371843 420639 371849
rect 420547 371809 420559 371843
rect 420627 371809 420639 371843
rect 420547 371803 420639 371809
rect 420394 371771 420426 371790
rect 420208 371759 420261 371771
rect 420208 371699 420221 371759
rect 420255 371699 420261 371759
rect 420208 371687 420261 371699
rect 420373 371759 420426 371771
rect 420373 371699 420379 371759
rect 420413 371699 420426 371759
rect 420373 371687 420426 371699
rect 420208 371660 420238 371687
rect 420000 371655 420080 371656
rect 419995 371649 420087 371655
rect 419995 371615 420007 371649
rect 420075 371642 420087 371649
rect 419995 371609 420008 371615
rect 420000 371586 420008 371609
rect 420076 371609 420087 371642
rect 420271 371649 420363 371655
rect 420271 371615 420283 371649
rect 420351 371615 420363 371649
rect 420271 371609 420363 371615
rect 420076 371586 420080 371609
rect 420000 371578 420080 371586
rect 420394 371434 420426 371687
rect 420482 371771 420514 371788
rect 420668 371771 420698 371996
rect 420482 371759 420537 371771
rect 420482 371699 420497 371759
rect 420531 371699 420537 371759
rect 420482 371687 420537 371699
rect 420649 371759 420698 371771
rect 420649 371699 420655 371759
rect 420689 371699 420698 371759
rect 420649 371687 420698 371699
rect 420482 371434 420514 371687
rect 420668 371672 420698 371687
rect 420758 371771 420788 371996
rect 420823 371843 420915 371849
rect 420823 371809 420835 371843
rect 420903 371809 420915 371843
rect 420823 371803 420915 371809
rect 421099 371843 421191 371849
rect 421099 371809 421111 371843
rect 421179 371809 421191 371843
rect 421099 371803 421191 371809
rect 420946 371771 420978 371790
rect 420758 371759 420813 371771
rect 420758 371699 420773 371759
rect 420807 371699 420813 371759
rect 420758 371687 420813 371699
rect 420925 371759 420978 371771
rect 420925 371699 420931 371759
rect 420965 371699 420978 371759
rect 420925 371687 420978 371699
rect 420758 371672 420788 371687
rect 420547 371649 420639 371655
rect 420547 371615 420559 371649
rect 420627 371615 420639 371649
rect 420547 371609 420639 371615
rect 420823 371649 420915 371655
rect 420823 371615 420835 371649
rect 420903 371615 420915 371649
rect 420823 371609 420915 371615
rect 420946 371434 420978 371687
rect 421030 371771 421062 371782
rect 421222 371771 421252 371996
rect 421030 371759 421089 371771
rect 421030 371699 421049 371759
rect 421083 371699 421089 371759
rect 421030 371687 421089 371699
rect 421201 371759 421252 371771
rect 421201 371699 421207 371759
rect 421241 371699 421252 371759
rect 421201 371687 421252 371699
rect 421030 371434 421062 371687
rect 421222 371672 421252 371687
rect 421306 371771 421336 371996
rect 421375 371843 421467 371849
rect 421375 371809 421387 371843
rect 421455 371809 421467 371843
rect 421375 371803 421467 371809
rect 421496 371771 421528 371790
rect 421306 371759 421365 371771
rect 421306 371699 421325 371759
rect 421359 371699 421365 371759
rect 421306 371687 421365 371699
rect 421477 371759 421528 371771
rect 421477 371699 421483 371759
rect 421517 371699 421528 371759
rect 421477 371687 421528 371699
rect 421306 371674 421336 371687
rect 421099 371649 421191 371655
rect 421099 371615 421111 371649
rect 421179 371615 421191 371649
rect 421099 371609 421191 371615
rect 421375 371649 421467 371655
rect 421375 371615 421387 371649
rect 421455 371615 421467 371649
rect 421375 371609 421467 371615
rect 421496 371434 421528 371687
rect 421620 371576 421658 371996
rect 422747 371818 422801 371996
rect 508118 371900 508178 372060
rect 508338 371900 508924 372060
rect 509380 372016 509564 373280
rect 510030 372060 510570 372100
rect 509380 371924 509573 372016
rect 508118 371860 508924 371900
rect 508478 371854 508924 371860
rect 422668 371786 422868 371818
rect 508723 371816 508923 371854
rect 509395 371844 509573 371924
rect 422668 371638 422696 371786
rect 422844 371638 422868 371786
rect 422668 371618 422868 371638
rect 508821 371610 508851 371816
rect 509395 371784 509441 371844
rect 509535 371784 509573 371844
rect 510030 371900 510378 372060
rect 510538 371900 510570 372060
rect 510030 371842 510570 371900
rect 510073 371816 510273 371842
rect 509395 371750 509573 371784
rect 508821 371582 509971 371610
rect 508821 371443 508851 371582
rect 508890 371515 508982 371521
rect 508890 371481 508902 371515
rect 508970 371481 508982 371515
rect 508890 371475 508982 371481
rect 509166 371515 509258 371521
rect 509166 371481 509178 371515
rect 509246 371481 509258 371515
rect 509166 371475 509258 371481
rect 509015 371443 509049 371446
rect 418039 371388 421532 371434
rect 508821 371431 508880 371443
rect 421030 371386 421062 371388
rect 508821 371371 508840 371431
rect 508874 371371 508880 371431
rect 508821 371368 508880 371371
rect 338790 371278 339590 371364
rect 508834 371359 508880 371368
rect 508992 371431 509049 371443
rect 508992 371371 508998 371431
rect 509032 371412 509049 371431
rect 509101 371443 509137 371448
rect 509293 371443 509327 371582
rect 509101 371431 509156 371443
rect 509032 371371 509051 371412
rect 508992 371359 509051 371371
rect 419538 371334 419660 371344
rect 419538 371290 419566 371334
rect 419638 371290 419660 371334
rect 419538 371108 419660 371290
rect 508890 371321 508982 371327
rect 508890 371287 508902 371321
rect 508970 371287 508982 371321
rect 420000 371270 420090 371286
rect 508890 371281 508982 371287
rect 420000 371206 420012 371270
rect 420084 371206 420090 371270
rect 419504 371100 419704 371108
rect 232698 370957 232790 370963
rect 232698 370923 232710 370957
rect 232778 370923 232790 370957
rect 232698 370917 232790 370923
rect 232823 370885 232863 371061
rect 232642 370873 232688 370885
rect 230433 370815 232648 370873
rect 230433 370798 231381 370815
rect 141258 368634 142348 368640
rect 143138 370215 147492 370415
rect 143138 365815 143338 370215
rect 232484 370637 232526 370815
rect 232642 370813 232648 370815
rect 232682 370813 232688 370873
rect 232642 370801 232688 370813
rect 232800 370873 232863 370885
rect 232800 370813 232806 370873
rect 232840 370813 232863 370873
rect 232800 370801 232863 370813
rect 232823 370795 232863 370801
rect 232905 370885 232945 371061
rect 232974 370957 233066 370963
rect 232974 370923 232986 370957
rect 233054 370923 233066 370957
rect 232974 370917 233066 370923
rect 233250 370957 233342 370963
rect 233250 370923 233262 370957
rect 233330 370923 233342 370957
rect 233250 370917 233342 370923
rect 233099 370885 233129 370893
rect 232905 370873 232964 370885
rect 232905 370813 232924 370873
rect 232958 370813 232964 370873
rect 232905 370801 232964 370813
rect 233076 370873 233129 370885
rect 233076 370813 233082 370873
rect 233116 370813 233129 370873
rect 233076 370801 233129 370813
rect 232905 370797 232945 370801
rect 232698 370763 232790 370769
rect 232698 370729 232710 370763
rect 232778 370729 232790 370763
rect 232698 370723 232790 370729
rect 232974 370763 233066 370769
rect 232974 370729 232986 370763
rect 233054 370729 233066 370763
rect 232974 370723 233066 370729
rect 233099 370637 233129 370801
rect 233185 370885 233215 370893
rect 233381 370885 233421 371061
rect 233185 370873 233240 370885
rect 233185 370813 233200 370873
rect 233234 370813 233240 370873
rect 233185 370801 233240 370813
rect 233352 370873 233421 370885
rect 233352 370813 233358 370873
rect 233392 370813 233421 370873
rect 233352 370801 233421 370813
rect 233185 370637 233215 370801
rect 233381 370797 233421 370801
rect 233449 370885 233489 371061
rect 233526 370957 233618 370963
rect 233526 370923 233538 370957
rect 233606 370923 233618 370957
rect 233526 370917 233618 370923
rect 233802 370957 233894 370963
rect 233802 370923 233814 370957
rect 233882 370923 233894 370957
rect 233802 370917 233894 370923
rect 233653 370885 233683 370893
rect 233449 370873 233516 370885
rect 233449 370813 233476 370873
rect 233510 370813 233516 370873
rect 233449 370801 233516 370813
rect 233628 370873 233683 370885
rect 233628 370813 233634 370873
rect 233668 370813 233683 370873
rect 233628 370801 233683 370813
rect 233449 370797 233489 370801
rect 233250 370763 233342 370769
rect 233250 370729 233262 370763
rect 233330 370729 233342 370763
rect 233250 370723 233342 370729
rect 233526 370763 233618 370769
rect 233526 370729 233538 370763
rect 233606 370729 233618 370763
rect 233526 370723 233618 370729
rect 233653 370637 233683 370801
rect 233739 370885 233769 370893
rect 233929 370885 233969 371061
rect 233739 370873 233792 370885
rect 233739 370813 233752 370873
rect 233786 370813 233792 370873
rect 233739 370801 233792 370813
rect 233904 370873 233969 370885
rect 233904 370813 233910 370873
rect 233944 370813 233969 370873
rect 233904 370801 233969 370813
rect 233739 370637 233769 370801
rect 233929 370793 233969 370801
rect 234001 370885 234041 371061
rect 234078 370957 234170 370963
rect 234078 370923 234090 370957
rect 234158 370923 234170 370957
rect 234078 370917 234170 370923
rect 234354 370957 234446 370963
rect 234354 370923 234366 370957
rect 234434 370923 234446 370957
rect 234354 370917 234446 370923
rect 234201 370885 234231 370893
rect 234001 370873 234068 370885
rect 234001 370813 234028 370873
rect 234062 370813 234068 370873
rect 234001 370801 234068 370813
rect 234180 370873 234231 370885
rect 234180 370813 234186 370873
rect 234220 370813 234231 370873
rect 234180 370801 234231 370813
rect 234001 370797 234041 370801
rect 233802 370763 233894 370769
rect 233802 370729 233814 370763
rect 233882 370729 233894 370763
rect 233802 370723 233894 370729
rect 234078 370763 234170 370769
rect 234078 370729 234090 370763
rect 234158 370729 234170 370763
rect 234078 370723 234170 370729
rect 234201 370637 234231 370801
rect 234293 370885 234323 370891
rect 234481 370885 234521 371061
rect 234293 370873 234344 370885
rect 234293 370813 234304 370873
rect 234338 370813 234344 370873
rect 234293 370801 234344 370813
rect 234456 370873 234521 370885
rect 234456 370813 234462 370873
rect 234496 370813 234521 370873
rect 234456 370801 234521 370813
rect 234561 370885 234601 371061
rect 234630 370957 234722 370963
rect 234630 370923 234642 370957
rect 234710 370923 234722 370957
rect 234630 370917 234722 370923
rect 234906 370957 234998 370963
rect 234906 370923 234918 370957
rect 234986 370923 234998 370957
rect 234906 370917 234998 370923
rect 234751 370885 234781 370891
rect 234561 370873 234620 370885
rect 234561 370813 234580 370873
rect 234614 370813 234620 370873
rect 234561 370801 234620 370813
rect 234732 370873 234781 370885
rect 234732 370813 234738 370873
rect 234772 370813 234781 370873
rect 234732 370801 234781 370813
rect 234293 370637 234323 370801
rect 234354 370763 234446 370769
rect 234354 370729 234366 370763
rect 234434 370729 234446 370763
rect 234354 370723 234446 370729
rect 234630 370763 234722 370769
rect 234630 370729 234642 370763
rect 234710 370729 234722 370763
rect 234630 370723 234722 370729
rect 234751 370637 234781 370801
rect 234843 370885 234873 370889
rect 235035 370885 235075 371061
rect 234843 370873 234896 370885
rect 234843 370813 234856 370873
rect 234890 370813 234896 370873
rect 234843 370801 234896 370813
rect 235008 370873 235075 370885
rect 235008 370813 235014 370873
rect 235048 370813 235075 370873
rect 235008 370801 235075 370813
rect 234843 370637 234873 370801
rect 235035 370797 235075 370801
rect 235109 370885 235149 371061
rect 235182 370957 235274 370963
rect 235182 370923 235194 370957
rect 235262 370923 235274 370957
rect 235182 370917 235274 370923
rect 235458 370957 235550 370963
rect 235458 370923 235470 370957
rect 235538 370923 235550 370957
rect 235458 370917 235550 370923
rect 235307 370885 235337 370889
rect 235109 370873 235172 370885
rect 235109 370813 235132 370873
rect 235166 370813 235172 370873
rect 235109 370801 235172 370813
rect 235284 370873 235337 370885
rect 235284 370813 235290 370873
rect 235324 370813 235337 370873
rect 235284 370801 235337 370813
rect 235109 370799 235149 370801
rect 234906 370763 234998 370769
rect 234906 370729 234918 370763
rect 234986 370729 234998 370763
rect 234906 370723 234998 370729
rect 235182 370763 235274 370769
rect 235182 370729 235194 370763
rect 235262 370729 235274 370763
rect 235182 370723 235274 370729
rect 235307 370637 235337 370801
rect 235395 370885 235425 370887
rect 235587 370885 235627 371061
rect 235395 370873 235448 370885
rect 235395 370813 235408 370873
rect 235442 370813 235448 370873
rect 235395 370801 235448 370813
rect 235560 370873 235627 370885
rect 235560 370813 235566 370873
rect 235600 370813 235627 370873
rect 235560 370801 235627 370813
rect 235395 370637 235425 370801
rect 235587 370795 235627 370801
rect 235657 370885 235697 371061
rect 235734 370957 235826 370963
rect 235734 370923 235746 370957
rect 235814 370923 235826 370957
rect 235734 370917 235826 370923
rect 236010 370957 236102 370963
rect 236010 370923 236022 370957
rect 236090 370923 236102 370957
rect 236010 370917 236102 370923
rect 235857 370885 235887 370887
rect 235657 370873 235724 370885
rect 235657 370813 235684 370873
rect 235718 370813 235724 370873
rect 235657 370801 235724 370813
rect 235836 370873 235887 370885
rect 235836 370813 235842 370873
rect 235876 370813 235887 370873
rect 235836 370801 235887 370813
rect 235657 370799 235697 370801
rect 235458 370763 235550 370769
rect 235734 370767 235826 370769
rect 235458 370729 235470 370763
rect 235538 370729 235550 370763
rect 235731 370763 235826 370767
rect 235731 370734 235746 370763
rect 235458 370723 235550 370729
rect 235734 370729 235746 370734
rect 235814 370729 235826 370763
rect 235734 370723 235826 370729
rect 235857 370637 235887 370801
rect 235945 370885 235975 370887
rect 236135 370885 236175 371061
rect 235945 370873 236000 370885
rect 235945 370813 235960 370873
rect 235994 370813 236000 370873
rect 235945 370801 236000 370813
rect 236112 370873 236175 370885
rect 236112 370813 236118 370873
rect 236152 370813 236175 370873
rect 236112 370801 236175 370813
rect 235945 370637 235975 370801
rect 236135 370795 236175 370801
rect 236213 370885 236253 371061
rect 236286 370957 236378 370963
rect 236286 370923 236298 370957
rect 236366 370923 236378 370957
rect 236286 370917 236378 370923
rect 236562 370957 236654 370963
rect 236562 370923 236574 370957
rect 236642 370923 236654 370957
rect 236562 370917 236654 370923
rect 236409 370885 236439 370889
rect 236213 370873 236276 370885
rect 236213 370813 236236 370873
rect 236270 370813 236276 370873
rect 236213 370801 236276 370813
rect 236388 370873 236439 370885
rect 236388 370813 236394 370873
rect 236428 370813 236439 370873
rect 236388 370801 236439 370813
rect 236213 370799 236253 370801
rect 236010 370763 236102 370769
rect 236010 370729 236022 370763
rect 236090 370729 236102 370763
rect 236010 370723 236102 370729
rect 236286 370763 236378 370769
rect 236286 370729 236298 370763
rect 236366 370729 236378 370763
rect 236286 370723 236378 370729
rect 236409 370637 236439 370801
rect 236497 370885 236527 370889
rect 236689 370885 236729 371061
rect 236497 370873 236552 370885
rect 236497 370813 236512 370873
rect 236546 370813 236552 370873
rect 236497 370801 236552 370813
rect 236664 370873 236729 370885
rect 236664 370813 236670 370873
rect 236704 370813 236729 370873
rect 236664 370801 236729 370813
rect 236497 370637 236527 370801
rect 236689 370787 236729 370801
rect 236767 370885 236807 371061
rect 236838 370957 236930 370963
rect 236838 370923 236850 370957
rect 236918 370923 236930 370957
rect 236838 370917 236930 370923
rect 237114 370957 237206 370963
rect 237114 370923 237126 370957
rect 237194 370923 237206 370957
rect 237114 370917 237206 370923
rect 236961 370885 236991 370889
rect 236767 370873 236828 370885
rect 236767 370813 236788 370873
rect 236822 370813 236828 370873
rect 236767 370801 236828 370813
rect 236940 370873 236991 370885
rect 236940 370813 236946 370873
rect 236980 370813 236991 370873
rect 236940 370801 236991 370813
rect 236767 370795 236807 370801
rect 236562 370763 236654 370769
rect 236562 370729 236574 370763
rect 236642 370729 236654 370763
rect 236562 370723 236654 370729
rect 236838 370763 236930 370769
rect 236838 370729 236850 370763
rect 236918 370729 236930 370763
rect 236838 370723 236930 370729
rect 236961 370637 236991 370801
rect 237053 370885 237083 370889
rect 237245 370885 237285 371061
rect 237053 370873 237104 370885
rect 237053 370813 237064 370873
rect 237098 370813 237104 370873
rect 237053 370801 237104 370813
rect 237216 370873 237285 370885
rect 237216 370813 237222 370873
rect 237256 370813 237285 370873
rect 237216 370801 237285 370813
rect 237319 370885 237359 371061
rect 237390 370957 237482 370963
rect 237390 370923 237402 370957
rect 237470 370923 237482 370957
rect 237390 370917 237482 370923
rect 237666 370957 237758 370963
rect 237666 370923 237678 370957
rect 237746 370923 237758 370957
rect 237666 370917 237758 370923
rect 237515 370885 237545 370899
rect 237319 370873 237380 370885
rect 237319 370813 237340 370873
rect 237374 370813 237380 370873
rect 237319 370801 237380 370813
rect 237492 370873 237545 370885
rect 237492 370813 237498 370873
rect 237532 370813 237545 370873
rect 237492 370801 237545 370813
rect 237053 370637 237083 370801
rect 237245 370797 237285 370801
rect 237114 370763 237206 370769
rect 237114 370729 237126 370763
rect 237194 370729 237206 370763
rect 237114 370723 237206 370729
rect 237390 370763 237482 370769
rect 237390 370729 237402 370763
rect 237470 370729 237482 370763
rect 237390 370723 237482 370729
rect 237515 370637 237545 370801
rect 237601 370885 237631 370897
rect 237789 370885 237823 371061
rect 237601 370873 237656 370885
rect 237601 370813 237616 370873
rect 237650 370813 237656 370873
rect 237601 370801 237656 370813
rect 237768 370873 237823 370885
rect 237768 370813 237774 370873
rect 237808 370813 237823 370873
rect 237768 370801 237823 370813
rect 237601 370637 237631 370801
rect 237789 370797 237823 370801
rect 237879 370885 237913 371061
rect 237942 370957 238034 370963
rect 237942 370923 237954 370957
rect 238022 370923 238034 370957
rect 237942 370917 238034 370923
rect 238218 370957 238310 370963
rect 238218 370923 238230 370957
rect 238298 370923 238310 370957
rect 238218 370917 238310 370923
rect 238069 370885 238099 370895
rect 237879 370873 237932 370885
rect 237879 370813 237892 370873
rect 237926 370813 237932 370873
rect 237879 370801 237932 370813
rect 238044 370873 238099 370885
rect 238044 370813 238050 370873
rect 238084 370813 238099 370873
rect 238044 370801 238099 370813
rect 237879 370797 237913 370801
rect 237666 370763 237758 370769
rect 237666 370729 237678 370763
rect 237746 370729 237758 370763
rect 237666 370723 237758 370729
rect 237942 370763 238034 370769
rect 237942 370729 237954 370763
rect 238022 370729 238034 370763
rect 237942 370723 238034 370729
rect 238069 370637 238099 370801
rect 238155 370885 238185 370895
rect 238345 370885 238379 371061
rect 238155 370873 238208 370885
rect 238155 370813 238168 370873
rect 238202 370813 238208 370873
rect 238155 370801 238208 370813
rect 238320 370873 238379 370885
rect 238320 370813 238326 370873
rect 238360 370813 238379 370873
rect 238320 370801 238379 370813
rect 238429 370885 238463 371061
rect 238494 370957 238586 370963
rect 238494 370923 238506 370957
rect 238574 370923 238586 370957
rect 238494 370917 238586 370923
rect 238621 370885 238655 370899
rect 238429 370873 238484 370885
rect 238429 370813 238444 370873
rect 238478 370813 238484 370873
rect 238429 370801 238484 370813
rect 238596 370873 238655 370885
rect 238596 370813 238602 370873
rect 238636 370813 238655 370873
rect 238596 370801 238655 370813
rect 238155 370637 238185 370801
rect 238345 370797 238379 370801
rect 238218 370763 238310 370769
rect 238218 370729 238230 370763
rect 238298 370729 238310 370763
rect 238218 370723 238310 370729
rect 238494 370763 238586 370769
rect 238494 370729 238506 370763
rect 238574 370729 238586 370763
rect 238494 370723 238586 370729
rect 238621 370637 238655 370801
rect 238703 370885 238737 371061
rect 238770 370957 238862 370963
rect 238770 370923 238782 370957
rect 238850 370923 238862 370957
rect 238770 370917 238862 370923
rect 239046 370957 239138 370963
rect 239046 370923 239058 370957
rect 239126 370923 239138 370957
rect 239046 370917 239138 370923
rect 238895 370885 238925 370897
rect 238703 370873 238760 370885
rect 238703 370813 238720 370873
rect 238754 370813 238760 370873
rect 238703 370801 238760 370813
rect 238872 370873 238925 370885
rect 238872 370813 238878 370873
rect 238912 370813 238925 370873
rect 238872 370801 238925 370813
rect 238703 370799 238737 370801
rect 238770 370763 238862 370769
rect 238770 370729 238782 370763
rect 238850 370729 238862 370763
rect 238770 370723 238862 370729
rect 238895 370637 238925 370801
rect 238983 370885 239013 370899
rect 239173 370885 239207 371061
rect 238983 370873 239036 370885
rect 238983 370813 238996 370873
rect 239030 370813 239036 370873
rect 238983 370801 239036 370813
rect 239148 370873 239207 370885
rect 239148 370813 239154 370873
rect 239188 370813 239207 370873
rect 239148 370801 239207 370813
rect 239259 370885 239293 371061
rect 239331 370999 239546 371009
rect 239331 370963 239461 370999
rect 239322 370957 239461 370963
rect 239322 370923 239334 370957
rect 239402 370939 239461 370957
rect 239521 370939 239546 370999
rect 239402 370929 239546 370939
rect 239598 370957 239690 370963
rect 239402 370923 239414 370929
rect 239322 370917 239414 370923
rect 239598 370923 239610 370957
rect 239678 370923 239690 370957
rect 239598 370917 239690 370923
rect 239443 370885 239473 370899
rect 239259 370873 239312 370885
rect 239259 370813 239272 370873
rect 239306 370813 239312 370873
rect 239259 370801 239312 370813
rect 239424 370873 239473 370885
rect 239424 370813 239430 370873
rect 239464 370813 239473 370873
rect 239424 370801 239473 370813
rect 238983 370637 239013 370801
rect 239259 370795 239293 370801
rect 239046 370763 239138 370769
rect 239046 370729 239058 370763
rect 239126 370729 239138 370763
rect 239322 370763 239414 370769
rect 239322 370744 239334 370763
rect 239046 370723 239138 370729
rect 239186 370739 239334 370744
rect 239186 370684 239196 370739
rect 239261 370729 239334 370739
rect 239402 370729 239414 370763
rect 239261 370723 239414 370729
rect 239261 370694 239401 370723
rect 239261 370684 239271 370694
rect 239186 370679 239271 370684
rect 239443 370637 239473 370801
rect 239535 370885 239565 370899
rect 239725 370885 239759 371061
rect 239535 370873 239588 370885
rect 239535 370813 239548 370873
rect 239582 370813 239588 370873
rect 239535 370801 239588 370813
rect 239700 370873 239759 370885
rect 239700 370813 239706 370873
rect 239740 370813 239759 370873
rect 239700 370803 239759 370813
rect 239811 370885 239845 371061
rect 239874 370957 239966 370963
rect 239874 370923 239886 370957
rect 239954 370923 239966 370957
rect 239874 370917 239966 370923
rect 240150 370957 240242 370963
rect 240150 370923 240162 370957
rect 240230 370923 240242 370957
rect 240150 370917 240242 370923
rect 239997 370885 240027 370899
rect 239811 370873 239864 370885
rect 239811 370813 239824 370873
rect 239858 370813 239864 370873
rect 239700 370801 239746 370803
rect 239811 370801 239864 370813
rect 239976 370873 240027 370885
rect 239976 370813 239982 370873
rect 240016 370813 240027 370873
rect 239976 370801 240027 370813
rect 239535 370637 239565 370801
rect 239811 370799 239845 370801
rect 239598 370763 239690 370769
rect 239598 370729 239610 370763
rect 239678 370729 239690 370763
rect 239598 370723 239690 370729
rect 239874 370763 239966 370769
rect 239874 370729 239886 370763
rect 239954 370729 239966 370763
rect 239874 370723 239966 370729
rect 239997 370637 240027 370801
rect 240089 370885 240119 370899
rect 240275 370885 240309 371061
rect 240089 370873 240140 370885
rect 240089 370813 240100 370873
rect 240134 370813 240140 370873
rect 240089 370801 240140 370813
rect 240252 370873 240309 370885
rect 240252 370813 240258 370873
rect 240292 370813 240309 370873
rect 240252 370801 240309 370813
rect 240089 370637 240119 370801
rect 240275 370799 240309 370801
rect 240363 370885 240397 371061
rect 240426 370957 240518 370963
rect 240426 370923 240438 370957
rect 240506 370923 240518 370957
rect 240426 370917 240518 370923
rect 240702 370957 240794 370963
rect 240702 370923 240714 370957
rect 240782 370923 240794 370957
rect 240702 370917 240794 370923
rect 240549 370885 240579 370899
rect 240363 370873 240416 370885
rect 240363 370813 240376 370873
rect 240410 370813 240416 370873
rect 240363 370801 240416 370813
rect 240528 370873 240579 370885
rect 240528 370813 240534 370873
rect 240568 370813 240579 370873
rect 240528 370801 240579 370813
rect 240363 370797 240397 370801
rect 240150 370763 240242 370769
rect 240150 370729 240162 370763
rect 240230 370729 240242 370763
rect 240150 370723 240242 370729
rect 240426 370763 240518 370769
rect 240426 370729 240438 370763
rect 240506 370729 240518 370763
rect 240426 370723 240518 370729
rect 240549 370637 240579 370801
rect 240635 370885 240665 370899
rect 240831 370885 240865 371061
rect 240635 370873 240692 370885
rect 240635 370813 240652 370873
rect 240686 370813 240692 370873
rect 240635 370801 240692 370813
rect 240804 370873 240865 370885
rect 240804 370813 240810 370873
rect 240844 370813 240865 370873
rect 240804 370801 240865 370813
rect 240635 370637 240665 370801
rect 240831 370793 240865 370801
rect 240913 370885 240947 371061
rect 240978 370957 241070 370963
rect 240978 370923 240990 370957
rect 241058 370923 241070 370957
rect 240978 370917 241070 370923
rect 241254 370957 241346 370963
rect 241254 370923 241266 370957
rect 241334 370923 241346 370957
rect 241254 370917 241346 370923
rect 241103 370885 241133 370899
rect 240913 370873 240968 370885
rect 240913 370813 240928 370873
rect 240962 370813 240968 370873
rect 240913 370801 240968 370813
rect 241080 370873 241133 370885
rect 241080 370813 241086 370873
rect 241120 370813 241133 370873
rect 241080 370801 241133 370813
rect 240913 370799 240947 370801
rect 240702 370763 240794 370769
rect 240702 370729 240714 370763
rect 240782 370729 240794 370763
rect 240702 370723 240794 370729
rect 240978 370763 241070 370769
rect 240978 370729 240990 370763
rect 241058 370729 241070 370763
rect 240978 370723 241070 370729
rect 241103 370637 241133 370801
rect 241191 370885 241221 370897
rect 241385 370885 241419 371061
rect 241191 370873 241244 370885
rect 241191 370813 241204 370873
rect 241238 370813 241244 370873
rect 241191 370801 241244 370813
rect 241356 370873 241419 370885
rect 241356 370813 241362 370873
rect 241396 370813 241419 370873
rect 241356 370801 241419 370813
rect 241191 370637 241221 370801
rect 241385 370797 241419 370801
rect 241463 370885 241497 371061
rect 241530 370957 241622 370963
rect 241530 370923 241542 370957
rect 241610 370923 241622 370957
rect 241530 370917 241622 370923
rect 241806 370957 241898 370963
rect 241806 370923 241818 370957
rect 241886 370923 241898 370957
rect 241806 370917 241898 370923
rect 241655 370885 241685 370901
rect 241463 370873 241520 370885
rect 241463 370813 241480 370873
rect 241514 370813 241520 370873
rect 241463 370801 241520 370813
rect 241632 370873 241685 370885
rect 241632 370813 241638 370873
rect 241672 370813 241685 370873
rect 241632 370801 241685 370813
rect 241463 370799 241497 370801
rect 241254 370763 241346 370769
rect 241254 370729 241266 370763
rect 241334 370729 241346 370763
rect 241254 370723 241346 370729
rect 241530 370763 241622 370769
rect 241530 370729 241542 370763
rect 241610 370729 241622 370763
rect 241530 370723 241622 370729
rect 241655 370637 241685 370801
rect 241743 370885 241773 370901
rect 241941 370885 241975 371061
rect 241743 370873 241796 370885
rect 241743 370813 241756 370873
rect 241790 370813 241796 370873
rect 241743 370801 241796 370813
rect 241908 370873 241975 370885
rect 241908 370813 241914 370873
rect 241948 370813 241975 370873
rect 241908 370801 241975 370813
rect 241743 370637 241773 370801
rect 241941 370789 241975 370801
rect 242015 370885 242049 371061
rect 242082 370957 242174 370963
rect 242082 370923 242094 370957
rect 242162 370923 242174 370957
rect 242082 370917 242174 370923
rect 242358 370957 242450 370963
rect 242358 370923 242370 370957
rect 242438 370923 242450 370957
rect 242358 370917 242450 370923
rect 242205 370885 242235 370903
rect 242015 370873 242072 370885
rect 242015 370813 242032 370873
rect 242066 370813 242072 370873
rect 242015 370801 242072 370813
rect 242184 370873 242235 370885
rect 242184 370813 242190 370873
rect 242224 370813 242235 370873
rect 242184 370801 242235 370813
rect 242015 370793 242049 370801
rect 241806 370763 241898 370769
rect 241806 370729 241818 370763
rect 241886 370729 241898 370763
rect 241806 370723 241898 370729
rect 242082 370763 242174 370769
rect 242082 370729 242094 370763
rect 242162 370729 242174 370763
rect 242082 370723 242174 370729
rect 242205 370637 242235 370801
rect 242293 370885 242323 370901
rect 242485 370885 242519 371061
rect 242293 370873 242348 370885
rect 242293 370813 242308 370873
rect 242342 370813 242348 370873
rect 242293 370801 242348 370813
rect 242460 370873 242519 370885
rect 242460 370813 242466 370873
rect 242500 370813 242519 370873
rect 242460 370801 242519 370813
rect 242293 370637 242323 370801
rect 242485 370789 242519 370801
rect 242565 370885 242599 371061
rect 242634 370957 242726 370963
rect 242634 370923 242646 370957
rect 242714 370923 242726 370957
rect 242634 370917 242726 370923
rect 242910 370957 243002 370963
rect 242910 370923 242922 370957
rect 242990 370923 243002 370957
rect 242910 370917 243002 370923
rect 242757 370885 242787 370901
rect 242565 370873 242624 370885
rect 242565 370813 242584 370873
rect 242618 370813 242624 370873
rect 242565 370801 242624 370813
rect 242736 370873 242787 370885
rect 242736 370813 242742 370873
rect 242776 370813 242787 370873
rect 242736 370801 242787 370813
rect 242565 370787 242599 370801
rect 242358 370763 242450 370769
rect 242358 370729 242370 370763
rect 242438 370729 242450 370763
rect 242358 370723 242450 370729
rect 242634 370763 242726 370769
rect 242634 370729 242646 370763
rect 242714 370729 242726 370763
rect 242634 370723 242726 370729
rect 242757 370637 242787 370801
rect 242845 370885 242875 370903
rect 243041 370885 243075 371061
rect 242845 370873 242900 370885
rect 242845 370813 242860 370873
rect 242894 370813 242900 370873
rect 242845 370801 242900 370813
rect 243012 370873 243075 370885
rect 243012 370813 243018 370873
rect 243052 370813 243075 370873
rect 243012 370801 243075 370813
rect 242845 370637 242875 370801
rect 243041 370789 243075 370801
rect 243115 370885 243149 371061
rect 243186 370957 243278 370963
rect 243186 370923 243198 370957
rect 243266 370923 243278 370957
rect 243186 370917 243278 370923
rect 243462 370957 243554 370963
rect 243462 370923 243474 370957
rect 243542 370923 243554 370957
rect 243462 370917 243554 370923
rect 243309 370885 243339 370901
rect 243115 370873 243176 370885
rect 243115 370813 243136 370873
rect 243170 370813 243176 370873
rect 243115 370801 243176 370813
rect 243288 370873 243339 370885
rect 243288 370813 243294 370873
rect 243328 370813 243339 370873
rect 243288 370801 243339 370813
rect 243115 370787 243149 370801
rect 242910 370763 243002 370769
rect 242910 370729 242922 370763
rect 242990 370729 243002 370763
rect 242910 370723 243002 370729
rect 243186 370763 243278 370769
rect 243186 370729 243198 370763
rect 243266 370729 243278 370763
rect 243186 370723 243278 370729
rect 243309 370637 243339 370801
rect 243399 370885 243429 370903
rect 243591 370885 243625 371061
rect 243399 370873 243452 370885
rect 243399 370813 243412 370873
rect 243446 370813 243452 370873
rect 243399 370801 243452 370813
rect 243564 370873 243625 370885
rect 243564 370813 243570 370873
rect 243604 370813 243625 370873
rect 243564 370801 243625 370813
rect 243399 370637 243429 370801
rect 243591 370791 243625 370801
rect 243667 370885 243701 371061
rect 243738 370957 243830 370963
rect 243738 370923 243750 370957
rect 243818 370923 243830 370957
rect 243738 370917 243830 370923
rect 244014 370957 244106 370963
rect 244014 370923 244026 370957
rect 244094 370923 244106 370957
rect 244014 370917 244106 370923
rect 243861 370885 243891 370901
rect 243667 370873 243728 370885
rect 243667 370813 243688 370873
rect 243722 370813 243728 370873
rect 243667 370801 243728 370813
rect 243840 370873 243891 370885
rect 243840 370813 243846 370873
rect 243880 370813 243891 370873
rect 243840 370801 243891 370813
rect 243667 370791 243701 370801
rect 243462 370763 243554 370769
rect 243462 370729 243474 370763
rect 243542 370729 243554 370763
rect 243462 370723 243554 370729
rect 243738 370763 243830 370769
rect 243738 370729 243750 370763
rect 243818 370729 243830 370763
rect 243738 370723 243830 370729
rect 243861 370637 243891 370801
rect 243951 370885 243981 370903
rect 244141 370885 244175 371061
rect 243951 370873 244004 370885
rect 243951 370813 243964 370873
rect 243998 370813 244004 370873
rect 243951 370801 244004 370813
rect 244116 370873 244175 370885
rect 244116 370813 244122 370873
rect 244156 370813 244175 370873
rect 244116 370801 244175 370813
rect 243951 370637 243981 370801
rect 244141 370795 244175 370801
rect 244223 370885 244257 371061
rect 244290 370957 244382 370963
rect 244290 370923 244302 370957
rect 244370 370923 244382 370957
rect 244290 370917 244382 370923
rect 244566 370957 244658 370963
rect 244566 370923 244578 370957
rect 244646 370923 244658 370957
rect 244566 370917 244658 370923
rect 244415 370885 244445 370907
rect 244223 370873 244280 370885
rect 244223 370813 244240 370873
rect 244274 370813 244280 370873
rect 244223 370801 244280 370813
rect 244392 370873 244445 370885
rect 244392 370813 244398 370873
rect 244432 370813 244445 370873
rect 244392 370801 244445 370813
rect 244223 370793 244257 370801
rect 244014 370763 244106 370769
rect 244014 370729 244026 370763
rect 244094 370729 244106 370763
rect 244014 370723 244106 370729
rect 244290 370763 244382 370769
rect 244290 370729 244302 370763
rect 244370 370729 244382 370763
rect 244290 370723 244382 370729
rect 244415 370637 244445 370801
rect 244505 370885 244535 370909
rect 244693 370885 244727 371061
rect 244505 370873 244556 370885
rect 244505 370813 244516 370873
rect 244550 370813 244556 370873
rect 244505 370801 244556 370813
rect 244668 370873 244727 370885
rect 244668 370813 244674 370873
rect 244708 370813 244727 370873
rect 244668 370801 244727 370813
rect 244771 370885 244805 371061
rect 244842 370957 244934 370963
rect 244842 370923 244854 370957
rect 244922 370923 244934 370957
rect 244842 370917 244934 370923
rect 245118 370957 245210 370963
rect 245118 370923 245130 370957
rect 245198 370923 245210 370957
rect 245118 370917 245210 370923
rect 244969 370885 244999 370909
rect 244771 370873 244832 370885
rect 244771 370813 244792 370873
rect 244826 370813 244832 370873
rect 244771 370801 244832 370813
rect 244944 370873 244999 370885
rect 244944 370813 244950 370873
rect 244984 370813 244999 370873
rect 244944 370801 244999 370813
rect 244505 370637 244535 370801
rect 244693 370799 244727 370801
rect 244566 370763 244658 370769
rect 244566 370729 244578 370763
rect 244646 370729 244658 370763
rect 244566 370723 244658 370729
rect 244842 370763 244934 370769
rect 244842 370729 244854 370763
rect 244922 370729 244934 370763
rect 244842 370723 244934 370729
rect 244969 370637 244999 370801
rect 245055 370885 245085 370913
rect 245243 370885 245277 371061
rect 245055 370873 245108 370885
rect 245055 370813 245068 370873
rect 245102 370813 245108 370873
rect 245055 370801 245108 370813
rect 245220 370873 245277 370885
rect 245220 370813 245226 370873
rect 245260 370813 245277 370873
rect 245220 370801 245277 370813
rect 245055 370637 245085 370801
rect 245243 370797 245277 370801
rect 245327 370885 245361 371061
rect 245394 370957 245486 370963
rect 245394 370923 245406 370957
rect 245474 370923 245486 370957
rect 245394 370917 245486 370923
rect 245670 370957 245762 370963
rect 245670 370923 245682 370957
rect 245750 370923 245762 370957
rect 245670 370917 245762 370923
rect 245515 370885 245545 370899
rect 245327 370873 245384 370885
rect 245327 370813 245344 370873
rect 245378 370813 245384 370873
rect 245327 370801 245384 370813
rect 245496 370873 245545 370885
rect 245496 370813 245502 370873
rect 245536 370813 245545 370873
rect 245496 370801 245545 370813
rect 245327 370795 245361 370801
rect 245118 370763 245210 370769
rect 245118 370729 245130 370763
rect 245198 370729 245210 370763
rect 245118 370723 245210 370729
rect 245394 370763 245486 370769
rect 245394 370729 245406 370763
rect 245474 370729 245486 370763
rect 245394 370723 245486 370729
rect 245515 370637 245545 370801
rect 245607 370885 245637 370897
rect 245795 370885 245829 371061
rect 245607 370873 245660 370885
rect 245607 370813 245620 370873
rect 245654 370813 245660 370873
rect 245607 370801 245660 370813
rect 245772 370873 245829 370885
rect 245772 370813 245778 370873
rect 245812 370813 245829 370873
rect 245772 370801 245829 370813
rect 245607 370637 245637 370801
rect 245795 370797 245829 370801
rect 245879 370885 245913 371061
rect 245946 370957 246038 370963
rect 245946 370923 245958 370957
rect 246026 370923 246038 370957
rect 245946 370917 246038 370923
rect 246222 370957 246314 370963
rect 246222 370923 246234 370957
rect 246302 370923 246314 370957
rect 246222 370917 246314 370923
rect 246071 370885 246101 370899
rect 245879 370873 245936 370885
rect 245879 370813 245896 370873
rect 245930 370813 245936 370873
rect 245879 370801 245936 370813
rect 246048 370873 246101 370885
rect 246048 370813 246054 370873
rect 246088 370813 246101 370873
rect 246048 370801 246101 370813
rect 245879 370799 245913 370801
rect 245670 370763 245762 370769
rect 245670 370729 245682 370763
rect 245750 370729 245762 370763
rect 245670 370723 245762 370729
rect 245946 370763 246038 370769
rect 245946 370729 245958 370763
rect 246026 370729 246038 370763
rect 245946 370723 246038 370729
rect 246071 370637 246101 370801
rect 246155 370885 246185 370899
rect 246349 370885 246383 371061
rect 246155 370873 246212 370885
rect 246155 370813 246172 370873
rect 246206 370813 246212 370873
rect 246155 370801 246212 370813
rect 246324 370873 246383 370885
rect 246324 370813 246330 370873
rect 246364 370813 246383 370873
rect 246324 370803 246383 370813
rect 246427 370885 246461 371061
rect 246498 370957 246590 370963
rect 246498 370923 246510 370957
rect 246578 370923 246590 370957
rect 246498 370917 246590 370923
rect 246621 370885 246651 370899
rect 246427 370873 246488 370885
rect 246427 370813 246448 370873
rect 246482 370813 246488 370873
rect 246324 370801 246370 370803
rect 246427 370801 246488 370813
rect 246600 370873 246651 370885
rect 246600 370813 246606 370873
rect 246640 370813 246651 370873
rect 246600 370801 246651 370813
rect 246741 370809 246775 371061
rect 246155 370637 246185 370801
rect 246222 370763 246314 370769
rect 246222 370729 246234 370763
rect 246302 370729 246314 370763
rect 246222 370723 246314 370729
rect 246498 370763 246590 370769
rect 246498 370729 246510 370763
rect 246578 370729 246590 370763
rect 246498 370723 246590 370729
rect 246621 370637 246651 370801
rect 232484 370595 246653 370637
rect 246611 370593 246653 370595
rect 236663 370489 236803 370501
rect 236663 370433 236703 370489
rect 236781 370433 236803 370489
rect 236663 369819 236803 370433
rect 247591 370134 249092 371061
rect 158318 369724 159188 369730
rect 233035 369619 236849 369819
rect 233035 367388 233235 369619
rect 322870 370892 328032 371092
rect 418428 370908 419704 371100
rect 322870 369490 323194 370892
rect 418428 370882 419702 370908
rect 412872 370836 419702 370882
rect 412872 370618 418692 370836
rect 322872 369146 323136 369490
rect 412872 369146 413136 370618
rect 420000 370340 420090 371206
rect 508901 371244 508969 371281
rect 508901 371210 508923 371244
rect 508961 371210 508969 371244
rect 508901 371066 508969 371210
rect 509015 371175 509051 371359
rect 509101 371371 509116 371431
rect 509150 371371 509156 371431
rect 509101 371359 509156 371371
rect 509268 371431 509327 371443
rect 509268 371371 509274 371431
rect 509308 371371 509327 371431
rect 509268 371359 509327 371371
rect 509101 371175 509137 371359
rect 509293 371340 509327 371359
rect 509371 371443 509405 371582
rect 509437 371542 509539 371550
rect 509437 371484 509445 371542
rect 509531 371484 509539 371542
rect 509437 371481 509454 371484
rect 509522 371481 509539 371484
rect 509437 371476 509539 371481
rect 509718 371515 509810 371521
rect 509718 371481 509730 371515
rect 509798 371481 509810 371515
rect 509442 371475 509534 371476
rect 509718 371475 509810 371481
rect 509573 371443 509611 371444
rect 509851 371443 509885 371582
rect 509371 371431 509432 371443
rect 509371 371371 509392 371431
rect 509426 371371 509432 371431
rect 509371 371359 509432 371371
rect 509544 371431 509611 371443
rect 509662 371442 509708 371443
rect 509544 371371 509550 371431
rect 509584 371371 509611 371431
rect 509544 371359 509611 371371
rect 509371 371338 509405 371359
rect 509166 371321 509258 371327
rect 509442 371326 509534 371327
rect 509166 371287 509178 371321
rect 509246 371287 509258 371321
rect 509166 371281 509258 371287
rect 509437 371321 509539 371326
rect 509437 371318 509454 371321
rect 509522 371318 509539 371321
rect 509437 371260 509445 371318
rect 509531 371260 509539 371318
rect 509437 371252 509539 371260
rect 509015 371174 509295 371175
rect 509573 371174 509611 371359
rect 509647 371431 509708 371442
rect 509647 371371 509668 371431
rect 509702 371371 509708 371431
rect 509647 371359 509708 371371
rect 509820 371431 509885 371443
rect 509820 371371 509826 371431
rect 509860 371371 509885 371431
rect 509820 371359 509885 371371
rect 509647 371174 509685 371359
rect 509851 371340 509885 371359
rect 509921 371443 509955 371582
rect 509994 371515 510086 371521
rect 509994 371481 510006 371515
rect 510074 371481 510086 371515
rect 509994 371475 510086 371481
rect 510237 371444 510271 371816
rect 510117 371443 510271 371444
rect 509921 371431 509984 371443
rect 509921 371371 509944 371431
rect 509978 371371 509984 371431
rect 509921 371359 509984 371371
rect 510096 371434 510271 371443
rect 510096 371431 510269 371434
rect 510096 371371 510102 371431
rect 510136 371374 510269 371431
rect 510136 371371 510142 371374
rect 510096 371359 510142 371371
rect 509921 371344 509955 371359
rect 509718 371321 509810 371327
rect 509718 371287 509730 371321
rect 509798 371287 509810 371321
rect 509718 371281 509810 371287
rect 509994 371321 510086 371327
rect 509994 371287 510006 371321
rect 510074 371287 510086 371321
rect 509994 371281 510086 371287
rect 510237 371322 510269 371374
rect 510237 371174 510273 371322
rect 509015 371172 510273 371174
rect 509017 371142 510273 371172
rect 509017 371141 509585 371142
rect 509017 371138 509051 371141
rect 509293 371140 509585 371141
rect 508873 371044 509073 371066
rect 508812 370882 509076 371044
rect 509395 370996 509573 371026
rect 502872 370618 509076 370882
rect 509388 370990 509573 370996
rect 509388 370930 509439 370990
rect 509533 370930 509573 370990
rect 509388 370760 509573 370930
rect 417078 370336 419388 370340
rect 419652 370336 421758 370340
rect 417078 369740 421758 370336
rect 247591 368627 249092 368633
rect 52310 360230 53762 365815
rect 52310 359406 52640 360230
rect 53366 359406 53762 360230
rect 52310 358812 53762 359406
rect 142310 360230 143762 365815
rect 142310 359406 142640 360230
rect 143366 359406 143762 360230
rect 142310 358812 143762 359406
rect 232310 360230 233762 367388
rect 232310 359406 232640 360230
rect 233366 359406 233762 360230
rect 232310 358812 233762 359406
rect 322310 360230 323762 369146
rect 322310 359406 322640 360230
rect 323366 359406 323762 360230
rect 322310 358812 323762 359406
rect 412310 360230 413762 369146
rect 417078 368820 418038 369740
rect 417078 368220 417238 368820
rect 417838 368220 418038 368820
rect 417078 368060 418038 368220
rect 420798 368820 421758 369740
rect 502872 369146 503136 370618
rect 509388 370340 509564 370760
rect 507078 369740 511758 370340
rect 420798 368220 420958 368820
rect 421558 368220 421758 368820
rect 420798 368060 421758 368220
rect 412310 359406 412640 360230
rect 413366 359406 413762 360230
rect 412310 358812 413762 359406
rect 502310 360230 503762 369146
rect 507078 368820 508038 369740
rect 507078 368220 507238 368820
rect 507838 368220 508038 368820
rect 507078 368060 508038 368220
rect 510798 368820 511758 369740
rect 510798 368220 510958 368820
rect 511558 368220 511758 368820
rect 510798 368060 511758 368220
rect 502310 359406 502640 360230
rect 503366 359406 503762 360230
rect 502310 358812 503762 359406
rect 64394 264794 65846 265158
rect 64394 263970 64790 264794
rect 65516 263970 65846 264794
rect 57138 255400 58098 255560
rect 57138 254800 57298 255400
rect 57898 254800 58098 255400
rect 57138 253880 58098 254800
rect 60858 255400 61818 255560
rect 60858 254800 61018 255400
rect 61618 254800 61818 255400
rect 64394 254824 65846 263970
rect 153518 264590 154970 264954
rect 334394 264794 335846 265158
rect 153518 263766 153914 264590
rect 154640 263766 154970 264590
rect 146262 255196 147222 255356
rect 60858 253880 61818 254800
rect 57138 253280 61818 253880
rect 146262 254596 146422 255196
rect 147022 254596 147222 255196
rect 146262 253676 147222 254596
rect 149982 255196 150942 255356
rect 149982 254596 150142 255196
rect 150742 254596 150942 255196
rect 153518 254620 154970 263766
rect 244772 264402 246224 264766
rect 244772 263578 245168 264402
rect 245894 263578 246224 264402
rect 149982 253676 150942 254596
rect 244772 254432 246224 263578
rect 334394 263970 334790 264794
rect 335516 263970 335846 264794
rect 334394 255113 335846 263970
rect 424394 264794 425846 265158
rect 424394 263970 424790 264794
rect 425516 263970 425846 264794
rect 424394 258735 425846 263970
rect 514394 264794 515846 265158
rect 514394 263970 514790 264794
rect 515516 263970 515846 264794
rect 514394 258735 515846 263970
rect 58478 252100 58924 252104
rect 58118 252060 58924 252100
rect 58118 251900 58178 252060
rect 58338 251900 58924 252060
rect 59380 252016 59564 253280
rect 146262 253076 150942 253676
rect 234122 253110 234642 253344
rect 148504 252474 148688 253076
rect 234122 252986 234286 253110
rect 234394 252986 234642 253110
rect 148492 252388 149212 252474
rect 149126 252188 149212 252388
rect 234122 252308 234642 252986
rect 320433 252790 321381 252796
rect 149126 252124 149132 252188
rect 149204 252124 149212 252188
rect 234266 252206 234350 252308
rect 234266 252164 234282 252206
rect 234336 252164 234350 252206
rect 234266 252144 234350 252164
rect 60030 252060 60570 252100
rect 149126 252098 149212 252124
rect 59380 251924 59573 252016
rect 58118 251860 58924 251900
rect 58478 251854 58924 251860
rect 58723 251816 58923 251854
rect 59395 251844 59573 251924
rect 58821 251610 58851 251816
rect 59395 251784 59441 251844
rect 59535 251784 59573 251844
rect 60030 251900 60378 252060
rect 60538 251900 60570 252060
rect 249168 252008 249968 252142
rect 60030 251842 60570 251900
rect 60073 251816 60273 251842
rect 59395 251750 59573 251784
rect 58821 251582 59971 251610
rect 58821 251443 58851 251582
rect 58890 251515 58982 251521
rect 58890 251481 58902 251515
rect 58970 251481 58982 251515
rect 58890 251475 58982 251481
rect 59166 251515 59258 251521
rect 59166 251481 59178 251515
rect 59246 251481 59258 251515
rect 59166 251475 59258 251481
rect 59015 251443 59049 251446
rect 58821 251431 58880 251443
rect 58821 251371 58840 251431
rect 58874 251371 58880 251431
rect 58821 251368 58880 251371
rect 58834 251359 58880 251368
rect 58992 251431 59049 251443
rect 58992 251371 58998 251431
rect 59032 251412 59049 251431
rect 59101 251443 59137 251448
rect 59293 251443 59327 251582
rect 59101 251431 59156 251443
rect 59032 251371 59051 251412
rect 58992 251359 59051 251371
rect 58890 251321 58982 251327
rect 58890 251287 58902 251321
rect 58970 251287 58982 251321
rect 58890 251281 58982 251287
rect 58901 251244 58969 251281
rect 58901 251210 58923 251244
rect 58961 251210 58969 251244
rect 58901 251066 58969 251210
rect 59015 251175 59051 251359
rect 59101 251371 59116 251431
rect 59150 251371 59156 251431
rect 59101 251359 59156 251371
rect 59268 251431 59327 251443
rect 59268 251371 59274 251431
rect 59308 251371 59327 251431
rect 59268 251359 59327 251371
rect 59101 251175 59137 251359
rect 59293 251340 59327 251359
rect 59371 251443 59405 251582
rect 59437 251542 59539 251550
rect 59437 251484 59445 251542
rect 59531 251484 59539 251542
rect 59437 251481 59454 251484
rect 59522 251481 59539 251484
rect 59437 251476 59539 251481
rect 59718 251515 59810 251521
rect 59718 251481 59730 251515
rect 59798 251481 59810 251515
rect 59442 251475 59534 251476
rect 59718 251475 59810 251481
rect 59573 251443 59611 251444
rect 59851 251443 59885 251582
rect 59371 251431 59432 251443
rect 59371 251371 59392 251431
rect 59426 251371 59432 251431
rect 59371 251359 59432 251371
rect 59544 251431 59611 251443
rect 59662 251442 59708 251443
rect 59544 251371 59550 251431
rect 59584 251371 59611 251431
rect 59544 251359 59611 251371
rect 59371 251338 59405 251359
rect 59166 251321 59258 251327
rect 59442 251326 59534 251327
rect 59166 251287 59178 251321
rect 59246 251287 59258 251321
rect 59166 251281 59258 251287
rect 59437 251321 59539 251326
rect 59437 251318 59454 251321
rect 59522 251318 59539 251321
rect 59437 251260 59445 251318
rect 59531 251260 59539 251318
rect 59437 251252 59539 251260
rect 59015 251174 59295 251175
rect 59573 251174 59611 251359
rect 59647 251431 59708 251442
rect 59647 251371 59668 251431
rect 59702 251371 59708 251431
rect 59647 251359 59708 251371
rect 59820 251431 59885 251443
rect 59820 251371 59826 251431
rect 59860 251371 59885 251431
rect 59820 251359 59885 251371
rect 59647 251174 59685 251359
rect 59851 251340 59885 251359
rect 59921 251443 59955 251582
rect 59994 251515 60086 251521
rect 59994 251481 60006 251515
rect 60074 251481 60086 251515
rect 59994 251475 60086 251481
rect 60237 251444 60271 251816
rect 148130 251792 151928 251846
rect 148015 251639 148107 251645
rect 60117 251443 60271 251444
rect 59921 251431 59984 251443
rect 59921 251371 59944 251431
rect 59978 251371 59984 251431
rect 59921 251359 59984 251371
rect 60096 251434 60271 251443
rect 147088 251582 147288 251630
rect 148015 251605 148027 251639
rect 148095 251605 148107 251639
rect 148015 251599 148107 251605
rect 147088 251480 147120 251582
rect 147270 251480 147288 251582
rect 60096 251431 60269 251434
rect 60096 251371 60102 251431
rect 60136 251374 60269 251431
rect 147088 251430 147288 251480
rect 147952 251567 147984 251584
rect 148136 251567 148166 251792
rect 147952 251555 148005 251567
rect 147952 251495 147965 251555
rect 147999 251495 148005 251555
rect 147952 251483 148005 251495
rect 148117 251555 148166 251567
rect 148117 251495 148123 251555
rect 148157 251495 148166 251555
rect 148117 251483 148166 251495
rect 60136 251371 60142 251374
rect 60096 251359 60142 251371
rect 59921 251344 59955 251359
rect 59718 251321 59810 251327
rect 59718 251287 59730 251321
rect 59798 251287 59810 251321
rect 59718 251281 59810 251287
rect 59994 251321 60086 251327
rect 59994 251287 60006 251321
rect 60074 251287 60086 251321
rect 59994 251281 60086 251287
rect 60237 251322 60269 251374
rect 60237 251174 60273 251322
rect 147163 251230 147209 251430
rect 147952 251230 147984 251483
rect 148136 251462 148166 251483
rect 148226 251567 148256 251792
rect 148291 251639 148383 251645
rect 148291 251605 148303 251639
rect 148371 251605 148383 251639
rect 148291 251599 148383 251605
rect 148567 251639 148659 251645
rect 148567 251605 148579 251639
rect 148647 251605 148659 251639
rect 148567 251599 148659 251605
rect 148418 251567 148450 251586
rect 148226 251555 148281 251567
rect 148226 251495 148241 251555
rect 148275 251495 148281 251555
rect 148226 251483 148281 251495
rect 148393 251555 148450 251567
rect 148393 251495 148399 251555
rect 148433 251495 148450 251555
rect 148393 251483 148450 251495
rect 148226 251462 148256 251483
rect 148015 251445 148107 251451
rect 148015 251411 148027 251445
rect 148095 251411 148107 251445
rect 148015 251405 148107 251411
rect 148291 251445 148383 251451
rect 148291 251411 148303 251445
rect 148371 251411 148383 251445
rect 148291 251405 148383 251411
rect 148418 251230 148450 251483
rect 148500 251567 148532 251586
rect 148688 251567 148718 251792
rect 148500 251555 148557 251567
rect 148500 251495 148517 251555
rect 148551 251495 148557 251555
rect 148500 251483 148557 251495
rect 148669 251555 148718 251567
rect 148669 251495 148675 251555
rect 148709 251495 148718 251555
rect 148669 251483 148718 251495
rect 148500 251230 148532 251483
rect 148688 251464 148718 251483
rect 148778 251567 148808 251792
rect 149130 251668 149210 251678
rect 149130 251645 149132 251668
rect 148843 251639 148935 251645
rect 148843 251605 148855 251639
rect 148923 251605 148935 251639
rect 148843 251599 148935 251605
rect 149119 251639 149132 251645
rect 149200 251645 149210 251668
rect 149119 251605 149131 251639
rect 149200 251612 149211 251645
rect 149199 251605 149211 251612
rect 149119 251599 149211 251605
rect 148970 251567 149002 251586
rect 148778 251555 148833 251567
rect 148778 251495 148793 251555
rect 148827 251495 148833 251555
rect 148778 251483 148833 251495
rect 148945 251555 149002 251567
rect 148945 251495 148951 251555
rect 148985 251495 149002 251555
rect 148945 251483 149002 251495
rect 148778 251462 148808 251483
rect 148567 251445 148659 251451
rect 148567 251411 148579 251445
rect 148647 251411 148659 251445
rect 148567 251405 148659 251411
rect 148843 251445 148935 251451
rect 148843 251411 148855 251445
rect 148923 251411 148935 251445
rect 148843 251405 148935 251411
rect 148970 251230 149002 251483
rect 149058 251567 149090 251584
rect 149242 251567 149272 251792
rect 149058 251555 149109 251567
rect 149058 251495 149069 251555
rect 149103 251495 149109 251555
rect 149058 251483 149109 251495
rect 149221 251555 149272 251567
rect 149221 251495 149227 251555
rect 149261 251495 149272 251555
rect 149221 251483 149272 251495
rect 149058 251230 149090 251483
rect 149242 251458 149272 251483
rect 149332 251567 149362 251792
rect 149395 251639 149487 251645
rect 149395 251605 149407 251639
rect 149475 251605 149487 251639
rect 149395 251599 149487 251605
rect 149671 251639 149763 251645
rect 149671 251605 149683 251639
rect 149751 251605 149763 251639
rect 149671 251599 149763 251605
rect 149518 251567 149550 251586
rect 149332 251555 149385 251567
rect 149332 251495 149345 251555
rect 149379 251495 149385 251555
rect 149332 251483 149385 251495
rect 149497 251555 149550 251567
rect 149497 251495 149503 251555
rect 149537 251495 149550 251555
rect 149497 251483 149550 251495
rect 149332 251456 149362 251483
rect 149124 251451 149204 251452
rect 149119 251445 149211 251451
rect 149119 251411 149131 251445
rect 149199 251438 149211 251445
rect 149119 251405 149132 251411
rect 149124 251382 149132 251405
rect 149200 251405 149211 251438
rect 149395 251445 149487 251451
rect 149395 251411 149407 251445
rect 149475 251411 149487 251445
rect 149395 251405 149487 251411
rect 149200 251382 149204 251405
rect 149124 251374 149204 251382
rect 149518 251230 149550 251483
rect 149606 251567 149638 251584
rect 149792 251567 149822 251792
rect 149606 251555 149661 251567
rect 149606 251495 149621 251555
rect 149655 251495 149661 251555
rect 149606 251483 149661 251495
rect 149773 251555 149822 251567
rect 149773 251495 149779 251555
rect 149813 251495 149822 251555
rect 149773 251483 149822 251495
rect 149606 251230 149638 251483
rect 149792 251468 149822 251483
rect 149882 251567 149912 251792
rect 149947 251639 150039 251645
rect 149947 251605 149959 251639
rect 150027 251605 150039 251639
rect 149947 251599 150039 251605
rect 150223 251639 150315 251645
rect 150223 251605 150235 251639
rect 150303 251605 150315 251639
rect 150223 251599 150315 251605
rect 150070 251567 150102 251586
rect 149882 251555 149937 251567
rect 149882 251495 149897 251555
rect 149931 251495 149937 251555
rect 149882 251483 149937 251495
rect 150049 251555 150102 251567
rect 150049 251495 150055 251555
rect 150089 251495 150102 251555
rect 150049 251483 150102 251495
rect 149882 251468 149912 251483
rect 149671 251445 149763 251451
rect 149671 251411 149683 251445
rect 149751 251411 149763 251445
rect 149671 251405 149763 251411
rect 149947 251445 150039 251451
rect 149947 251411 149959 251445
rect 150027 251411 150039 251445
rect 149947 251405 150039 251411
rect 150070 251230 150102 251483
rect 150154 251567 150186 251578
rect 150346 251567 150376 251792
rect 150154 251555 150213 251567
rect 150154 251495 150173 251555
rect 150207 251495 150213 251555
rect 150154 251483 150213 251495
rect 150325 251555 150376 251567
rect 150325 251495 150331 251555
rect 150365 251495 150376 251555
rect 150325 251483 150376 251495
rect 150154 251230 150186 251483
rect 150346 251468 150376 251483
rect 150430 251567 150460 251792
rect 150499 251639 150591 251645
rect 150499 251605 150511 251639
rect 150579 251605 150591 251639
rect 150499 251599 150591 251605
rect 150620 251567 150652 251586
rect 150430 251555 150489 251567
rect 150430 251495 150449 251555
rect 150483 251495 150489 251555
rect 150430 251483 150489 251495
rect 150601 251555 150652 251567
rect 150601 251495 150607 251555
rect 150641 251495 150652 251555
rect 150601 251483 150652 251495
rect 150430 251470 150460 251483
rect 150223 251445 150315 251451
rect 150223 251411 150235 251445
rect 150303 251411 150315 251445
rect 150223 251405 150315 251411
rect 150499 251445 150591 251451
rect 150499 251411 150511 251445
rect 150579 251411 150591 251445
rect 150499 251405 150591 251411
rect 150620 251230 150652 251483
rect 150744 251372 150782 251792
rect 151871 251614 151925 251792
rect 232165 251636 232171 251962
rect 232497 251754 233034 251962
rect 234379 251942 249968 252008
rect 234259 251839 234351 251845
rect 234259 251805 234271 251839
rect 234339 251805 234351 251839
rect 234259 251799 234351 251805
rect 234384 251767 234424 251942
rect 234203 251755 234249 251767
rect 234203 251754 234209 251755
rect 232497 251696 234209 251754
rect 232497 251636 233034 251696
rect 151792 251582 151992 251614
rect 151792 251434 151820 251582
rect 151968 251434 151992 251582
rect 234045 251518 234087 251696
rect 234203 251695 234209 251696
rect 234243 251695 234249 251755
rect 234203 251683 234249 251695
rect 234361 251755 234424 251767
rect 234361 251695 234367 251755
rect 234401 251695 234424 251755
rect 234361 251683 234424 251695
rect 234384 251676 234424 251683
rect 234466 251767 234506 251942
rect 234535 251839 234627 251845
rect 234535 251805 234547 251839
rect 234615 251805 234627 251839
rect 234535 251799 234627 251805
rect 234811 251839 234903 251845
rect 234811 251805 234823 251839
rect 234891 251805 234903 251839
rect 234811 251799 234903 251805
rect 234660 251767 234690 251774
rect 234466 251755 234525 251767
rect 234466 251695 234485 251755
rect 234519 251695 234525 251755
rect 234466 251683 234525 251695
rect 234637 251755 234690 251767
rect 234637 251695 234643 251755
rect 234677 251695 234690 251755
rect 234637 251683 234690 251695
rect 234466 251678 234506 251683
rect 234259 251645 234351 251651
rect 234259 251611 234271 251645
rect 234339 251611 234351 251645
rect 234259 251605 234351 251611
rect 234535 251645 234627 251651
rect 234535 251611 234547 251645
rect 234615 251611 234627 251645
rect 234535 251605 234627 251611
rect 234217 251518 234393 251519
rect 234660 251518 234690 251683
rect 234746 251767 234776 251774
rect 234942 251767 234982 251942
rect 234746 251755 234801 251767
rect 234746 251695 234761 251755
rect 234795 251695 234801 251755
rect 234746 251683 234801 251695
rect 234913 251755 234982 251767
rect 234913 251695 234919 251755
rect 234953 251695 234982 251755
rect 234913 251683 234982 251695
rect 234746 251518 234776 251683
rect 234942 251678 234982 251683
rect 235010 251767 235050 251942
rect 235087 251839 235179 251845
rect 235087 251805 235099 251839
rect 235167 251805 235179 251839
rect 235087 251799 235179 251805
rect 235363 251839 235455 251845
rect 235363 251805 235375 251839
rect 235443 251805 235455 251839
rect 235363 251799 235455 251805
rect 235214 251767 235244 251774
rect 235010 251755 235077 251767
rect 235010 251695 235037 251755
rect 235071 251695 235077 251755
rect 235010 251683 235077 251695
rect 235189 251755 235244 251767
rect 235189 251695 235195 251755
rect 235229 251695 235244 251755
rect 235189 251683 235244 251695
rect 235010 251678 235050 251683
rect 234811 251645 234903 251651
rect 234811 251611 234823 251645
rect 234891 251611 234903 251645
rect 234811 251605 234903 251611
rect 235087 251645 235179 251651
rect 235087 251611 235099 251645
rect 235167 251611 235179 251645
rect 235087 251605 235179 251611
rect 235214 251518 235244 251683
rect 235300 251767 235330 251774
rect 235490 251767 235530 251942
rect 235300 251755 235353 251767
rect 235300 251695 235313 251755
rect 235347 251695 235353 251755
rect 235300 251683 235353 251695
rect 235465 251755 235530 251767
rect 235465 251695 235471 251755
rect 235505 251695 235530 251755
rect 235465 251683 235530 251695
rect 235300 251518 235330 251683
rect 235490 251674 235530 251683
rect 235562 251767 235602 251942
rect 235639 251839 235731 251845
rect 235639 251805 235651 251839
rect 235719 251805 235731 251839
rect 235639 251799 235731 251805
rect 235915 251839 236007 251845
rect 235915 251805 235927 251839
rect 235995 251805 236007 251839
rect 235915 251799 236007 251805
rect 235762 251767 235792 251774
rect 235562 251755 235629 251767
rect 235562 251695 235589 251755
rect 235623 251695 235629 251755
rect 235562 251683 235629 251695
rect 235741 251755 235792 251767
rect 235741 251695 235747 251755
rect 235781 251695 235792 251755
rect 235741 251683 235792 251695
rect 235562 251678 235602 251683
rect 235363 251645 235455 251651
rect 235363 251611 235375 251645
rect 235443 251611 235455 251645
rect 235363 251605 235455 251611
rect 235639 251645 235731 251651
rect 235639 251611 235651 251645
rect 235719 251611 235731 251645
rect 235639 251605 235731 251611
rect 235762 251518 235792 251683
rect 235854 251767 235884 251772
rect 236042 251767 236082 251942
rect 235854 251755 235905 251767
rect 235854 251695 235865 251755
rect 235899 251695 235905 251755
rect 235854 251683 235905 251695
rect 236017 251755 236082 251767
rect 236017 251695 236023 251755
rect 236057 251695 236082 251755
rect 236017 251683 236082 251695
rect 235854 251518 235884 251683
rect 236042 251682 236082 251683
rect 236122 251767 236162 251942
rect 236191 251839 236283 251845
rect 236191 251805 236203 251839
rect 236271 251805 236283 251839
rect 236191 251799 236283 251805
rect 236467 251839 236559 251845
rect 236467 251805 236479 251839
rect 236547 251805 236559 251839
rect 236467 251799 236559 251805
rect 236312 251767 236342 251772
rect 236122 251755 236181 251767
rect 236122 251695 236141 251755
rect 236175 251695 236181 251755
rect 236122 251683 236181 251695
rect 236293 251755 236342 251767
rect 236293 251695 236299 251755
rect 236333 251695 236342 251755
rect 236293 251683 236342 251695
rect 236122 251682 236162 251683
rect 235915 251645 236007 251651
rect 235915 251611 235927 251645
rect 235995 251611 236007 251645
rect 235915 251605 236007 251611
rect 236191 251645 236283 251651
rect 236191 251611 236203 251645
rect 236271 251611 236283 251645
rect 236191 251605 236283 251611
rect 236312 251518 236342 251683
rect 236404 251767 236434 251770
rect 236596 251767 236636 251942
rect 236404 251755 236457 251767
rect 236404 251695 236417 251755
rect 236451 251695 236457 251755
rect 236404 251683 236457 251695
rect 236569 251755 236636 251767
rect 236569 251695 236575 251755
rect 236609 251695 236636 251755
rect 236569 251683 236636 251695
rect 236404 251518 236434 251683
rect 236596 251678 236636 251683
rect 236670 251767 236710 251942
rect 236743 251839 236835 251845
rect 236743 251805 236755 251839
rect 236823 251805 236835 251839
rect 236743 251799 236835 251805
rect 237019 251839 237111 251845
rect 237019 251805 237031 251839
rect 237099 251805 237111 251839
rect 237019 251799 237111 251805
rect 236868 251767 236898 251770
rect 236670 251755 236733 251767
rect 236670 251695 236693 251755
rect 236727 251695 236733 251755
rect 236670 251683 236733 251695
rect 236845 251755 236898 251767
rect 236845 251695 236851 251755
rect 236885 251695 236898 251755
rect 236845 251683 236898 251695
rect 236670 251680 236710 251683
rect 236467 251645 236559 251651
rect 236467 251611 236479 251645
rect 236547 251611 236559 251645
rect 236467 251605 236559 251611
rect 236743 251645 236835 251651
rect 236743 251611 236755 251645
rect 236823 251611 236835 251645
rect 236743 251605 236835 251611
rect 236868 251518 236898 251683
rect 236956 251767 236986 251768
rect 237148 251767 237188 251942
rect 236956 251755 237009 251767
rect 236956 251695 236969 251755
rect 237003 251695 237009 251755
rect 236956 251683 237009 251695
rect 237121 251755 237188 251767
rect 237121 251695 237127 251755
rect 237161 251695 237188 251755
rect 237121 251683 237188 251695
rect 236956 251518 236986 251683
rect 237148 251676 237188 251683
rect 237218 251767 237258 251942
rect 237295 251839 237387 251845
rect 237295 251805 237307 251839
rect 237375 251805 237387 251839
rect 237295 251799 237387 251805
rect 237571 251839 237663 251845
rect 237571 251805 237583 251839
rect 237651 251805 237663 251839
rect 237571 251799 237663 251805
rect 237418 251767 237448 251768
rect 237218 251755 237285 251767
rect 237218 251695 237245 251755
rect 237279 251695 237285 251755
rect 237218 251683 237285 251695
rect 237397 251755 237448 251767
rect 237397 251695 237403 251755
rect 237437 251695 237448 251755
rect 237397 251683 237448 251695
rect 237218 251680 237258 251683
rect 237019 251645 237111 251651
rect 237019 251611 237031 251645
rect 237099 251611 237111 251645
rect 237019 251605 237111 251611
rect 237295 251645 237387 251651
rect 237295 251611 237307 251645
rect 237375 251611 237387 251645
rect 237295 251605 237387 251611
rect 237418 251518 237448 251683
rect 237506 251767 237536 251768
rect 237696 251767 237736 251942
rect 237506 251755 237561 251767
rect 237506 251695 237521 251755
rect 237555 251695 237561 251755
rect 237506 251683 237561 251695
rect 237673 251755 237736 251767
rect 237673 251695 237679 251755
rect 237713 251695 237736 251755
rect 237673 251683 237736 251695
rect 237506 251518 237536 251683
rect 237696 251676 237736 251683
rect 237774 251767 237814 251942
rect 237847 251839 237939 251845
rect 237847 251805 237859 251839
rect 237927 251805 237939 251839
rect 237847 251799 237939 251805
rect 238123 251839 238215 251845
rect 238123 251805 238135 251839
rect 238203 251805 238215 251839
rect 238123 251799 238215 251805
rect 237970 251767 238000 251770
rect 237774 251755 237837 251767
rect 237774 251695 237797 251755
rect 237831 251695 237837 251755
rect 237774 251683 237837 251695
rect 237949 251755 238000 251767
rect 237949 251695 237955 251755
rect 237989 251695 238000 251755
rect 237949 251683 238000 251695
rect 237774 251680 237814 251683
rect 237571 251645 237663 251651
rect 237571 251611 237583 251645
rect 237651 251611 237663 251645
rect 237571 251605 237663 251611
rect 237847 251645 237939 251651
rect 237847 251611 237859 251645
rect 237927 251611 237939 251645
rect 237847 251605 237939 251611
rect 237970 251518 238000 251683
rect 238058 251767 238088 251770
rect 238250 251767 238290 251942
rect 238058 251755 238113 251767
rect 238058 251695 238073 251755
rect 238107 251695 238113 251755
rect 238058 251683 238113 251695
rect 238225 251755 238290 251767
rect 238225 251695 238231 251755
rect 238265 251695 238290 251755
rect 238225 251683 238290 251695
rect 238058 251518 238088 251683
rect 238250 251668 238290 251683
rect 238328 251767 238368 251942
rect 238399 251839 238491 251845
rect 238399 251805 238411 251839
rect 238479 251805 238491 251839
rect 238399 251799 238491 251805
rect 238675 251839 238767 251845
rect 238675 251805 238687 251839
rect 238755 251805 238767 251839
rect 238675 251799 238767 251805
rect 238522 251767 238552 251770
rect 238328 251755 238389 251767
rect 238328 251695 238349 251755
rect 238383 251695 238389 251755
rect 238328 251683 238389 251695
rect 238501 251755 238552 251767
rect 238501 251695 238507 251755
rect 238541 251695 238552 251755
rect 238501 251683 238552 251695
rect 238328 251676 238368 251683
rect 238123 251645 238215 251651
rect 238123 251611 238135 251645
rect 238203 251611 238215 251645
rect 238123 251605 238215 251611
rect 238399 251645 238491 251651
rect 238399 251611 238411 251645
rect 238479 251611 238491 251645
rect 238399 251605 238491 251611
rect 238522 251518 238552 251683
rect 238614 251767 238644 251770
rect 238806 251767 238846 251942
rect 238614 251755 238665 251767
rect 238614 251695 238625 251755
rect 238659 251695 238665 251755
rect 238614 251683 238665 251695
rect 238777 251755 238846 251767
rect 238777 251695 238783 251755
rect 238817 251695 238846 251755
rect 238777 251683 238846 251695
rect 238614 251518 238644 251683
rect 238806 251678 238846 251683
rect 238880 251767 238920 251942
rect 238951 251839 239043 251845
rect 238951 251805 238963 251839
rect 239031 251805 239043 251839
rect 238951 251799 239043 251805
rect 239227 251839 239319 251845
rect 239227 251805 239239 251839
rect 239307 251805 239319 251839
rect 239227 251799 239319 251805
rect 239076 251767 239106 251780
rect 238880 251755 238941 251767
rect 238880 251695 238901 251755
rect 238935 251695 238941 251755
rect 238880 251683 238941 251695
rect 239053 251755 239106 251767
rect 239053 251695 239059 251755
rect 239093 251695 239106 251755
rect 239053 251683 239106 251695
rect 238880 251682 238920 251683
rect 238675 251645 238767 251651
rect 238675 251611 238687 251645
rect 238755 251611 238767 251645
rect 238675 251605 238767 251611
rect 238951 251645 239043 251651
rect 238951 251611 238963 251645
rect 239031 251611 239043 251645
rect 238951 251605 239043 251611
rect 239076 251518 239106 251683
rect 239162 251767 239192 251778
rect 239350 251767 239384 251942
rect 239162 251755 239217 251767
rect 239162 251695 239177 251755
rect 239211 251695 239217 251755
rect 239162 251683 239217 251695
rect 239329 251755 239384 251767
rect 239329 251695 239335 251755
rect 239369 251695 239384 251755
rect 239329 251683 239384 251695
rect 239162 251518 239192 251683
rect 239350 251678 239384 251683
rect 239440 251767 239474 251942
rect 239503 251839 239595 251845
rect 239503 251805 239515 251839
rect 239583 251805 239595 251839
rect 239503 251799 239595 251805
rect 239779 251839 239871 251845
rect 239779 251805 239791 251839
rect 239859 251805 239871 251839
rect 239779 251799 239871 251805
rect 239630 251767 239660 251776
rect 239440 251755 239493 251767
rect 239440 251695 239453 251755
rect 239487 251695 239493 251755
rect 239440 251683 239493 251695
rect 239605 251755 239660 251767
rect 239605 251695 239611 251755
rect 239645 251695 239660 251755
rect 239605 251683 239660 251695
rect 239440 251678 239474 251683
rect 239227 251645 239319 251651
rect 239227 251611 239239 251645
rect 239307 251611 239319 251645
rect 239227 251605 239319 251611
rect 239503 251645 239595 251651
rect 239503 251611 239515 251645
rect 239583 251611 239595 251645
rect 239503 251605 239595 251611
rect 239630 251518 239660 251683
rect 239716 251767 239746 251776
rect 239906 251767 239940 251942
rect 239716 251755 239769 251767
rect 239716 251695 239729 251755
rect 239763 251695 239769 251755
rect 239716 251683 239769 251695
rect 239881 251755 239940 251767
rect 239881 251695 239887 251755
rect 239921 251695 239940 251755
rect 239881 251683 239940 251695
rect 239716 251518 239746 251683
rect 239906 251678 239940 251683
rect 239990 251767 240024 251942
rect 240055 251839 240147 251845
rect 240055 251805 240067 251839
rect 240135 251805 240147 251839
rect 240055 251799 240147 251805
rect 240182 251767 240216 251780
rect 239990 251755 240045 251767
rect 239990 251695 240005 251755
rect 240039 251695 240045 251755
rect 239990 251683 240045 251695
rect 240157 251755 240216 251767
rect 240157 251695 240163 251755
rect 240197 251695 240216 251755
rect 240157 251683 240216 251695
rect 239990 251682 240024 251683
rect 239779 251645 239871 251651
rect 239779 251611 239791 251645
rect 239859 251611 239871 251645
rect 239779 251605 239871 251611
rect 240055 251645 240147 251651
rect 240055 251611 240067 251645
rect 240135 251611 240147 251645
rect 240055 251605 240147 251611
rect 240182 251518 240216 251683
rect 240264 251767 240298 251942
rect 240331 251839 240423 251845
rect 240331 251805 240343 251839
rect 240411 251805 240423 251839
rect 240331 251799 240423 251805
rect 240607 251839 240699 251845
rect 240607 251805 240619 251839
rect 240687 251805 240699 251839
rect 240607 251799 240699 251805
rect 240456 251767 240486 251778
rect 240264 251755 240321 251767
rect 240264 251695 240281 251755
rect 240315 251695 240321 251755
rect 240264 251683 240321 251695
rect 240433 251755 240486 251767
rect 240433 251695 240439 251755
rect 240473 251695 240486 251755
rect 240433 251683 240486 251695
rect 240264 251680 240298 251683
rect 240331 251645 240423 251651
rect 240331 251611 240343 251645
rect 240411 251611 240423 251645
rect 240331 251605 240423 251611
rect 240456 251518 240486 251683
rect 240544 251767 240574 251780
rect 240734 251767 240768 251942
rect 240544 251755 240597 251767
rect 240544 251695 240557 251755
rect 240591 251695 240597 251755
rect 240544 251683 240597 251695
rect 240709 251755 240768 251767
rect 240709 251695 240715 251755
rect 240749 251695 240768 251755
rect 240709 251683 240768 251695
rect 240544 251518 240574 251683
rect 240734 251682 240768 251683
rect 240820 251767 240854 251942
rect 240883 251839 240975 251845
rect 240883 251805 240895 251839
rect 240963 251805 240975 251839
rect 240883 251799 240975 251805
rect 241159 251839 241251 251845
rect 241159 251805 241171 251839
rect 241239 251805 241251 251839
rect 241159 251799 241251 251805
rect 241004 251767 241034 251780
rect 240820 251755 240873 251767
rect 240820 251695 240833 251755
rect 240867 251695 240873 251755
rect 240820 251683 240873 251695
rect 240985 251755 241034 251767
rect 240985 251695 240991 251755
rect 241025 251695 241034 251755
rect 240985 251683 241034 251695
rect 240820 251676 240854 251683
rect 240607 251645 240699 251651
rect 240607 251611 240619 251645
rect 240687 251611 240699 251645
rect 240607 251605 240699 251611
rect 240883 251645 240975 251651
rect 240883 251611 240895 251645
rect 240963 251611 240975 251645
rect 240883 251605 240975 251611
rect 241004 251518 241034 251683
rect 241096 251767 241126 251780
rect 241286 251767 241320 251942
rect 241096 251755 241149 251767
rect 241096 251695 241109 251755
rect 241143 251695 241149 251755
rect 241096 251683 241149 251695
rect 241261 251755 241320 251767
rect 241261 251695 241267 251755
rect 241301 251695 241320 251755
rect 241261 251684 241320 251695
rect 241372 251767 241406 251942
rect 241435 251839 241527 251845
rect 241435 251805 241447 251839
rect 241515 251805 241527 251839
rect 241435 251799 241527 251805
rect 241711 251839 241803 251845
rect 241711 251805 241723 251839
rect 241791 251805 241803 251839
rect 241711 251799 241803 251805
rect 241558 251767 241588 251780
rect 241372 251755 241425 251767
rect 241372 251695 241385 251755
rect 241419 251695 241425 251755
rect 241261 251683 241307 251684
rect 241372 251683 241425 251695
rect 241537 251755 241588 251767
rect 241537 251695 241543 251755
rect 241577 251695 241588 251755
rect 241537 251683 241588 251695
rect 241096 251518 241126 251683
rect 241372 251680 241406 251683
rect 241159 251645 241251 251651
rect 241159 251611 241171 251645
rect 241239 251611 241251 251645
rect 241159 251605 241251 251611
rect 241435 251645 241527 251651
rect 241435 251611 241447 251645
rect 241515 251611 241527 251645
rect 241435 251605 241527 251611
rect 241558 251518 241588 251683
rect 241650 251767 241680 251780
rect 241836 251767 241870 251942
rect 241650 251755 241701 251767
rect 241650 251695 241661 251755
rect 241695 251695 241701 251755
rect 241650 251683 241701 251695
rect 241813 251755 241870 251767
rect 241813 251695 241819 251755
rect 241853 251695 241870 251755
rect 241813 251683 241870 251695
rect 241650 251518 241680 251683
rect 241836 251680 241870 251683
rect 241924 251767 241958 251942
rect 241987 251839 242079 251845
rect 241987 251805 241999 251839
rect 242067 251805 242079 251839
rect 241987 251799 242079 251805
rect 242263 251839 242355 251845
rect 242263 251805 242275 251839
rect 242343 251805 242355 251839
rect 242263 251799 242355 251805
rect 242110 251767 242140 251780
rect 241924 251755 241977 251767
rect 241924 251695 241937 251755
rect 241971 251695 241977 251755
rect 241924 251683 241977 251695
rect 242089 251755 242140 251767
rect 242089 251695 242095 251755
rect 242129 251695 242140 251755
rect 242089 251683 242140 251695
rect 241924 251678 241958 251683
rect 241711 251645 241803 251651
rect 241711 251611 241723 251645
rect 241791 251611 241803 251645
rect 241711 251605 241803 251611
rect 241987 251645 242079 251651
rect 241987 251611 241999 251645
rect 242067 251611 242079 251645
rect 241987 251605 242079 251611
rect 242110 251518 242140 251683
rect 242196 251767 242226 251780
rect 242392 251767 242426 251942
rect 242196 251755 242253 251767
rect 242196 251695 242213 251755
rect 242247 251695 242253 251755
rect 242196 251683 242253 251695
rect 242365 251755 242426 251767
rect 242365 251695 242371 251755
rect 242405 251695 242426 251755
rect 242365 251683 242426 251695
rect 242196 251518 242226 251683
rect 242392 251674 242426 251683
rect 242474 251767 242508 251942
rect 242539 251839 242631 251845
rect 242539 251805 242551 251839
rect 242619 251805 242631 251839
rect 242539 251799 242631 251805
rect 242815 251839 242907 251845
rect 242815 251805 242827 251839
rect 242895 251805 242907 251839
rect 242815 251799 242907 251805
rect 242664 251767 242694 251780
rect 242474 251755 242529 251767
rect 242474 251695 242489 251755
rect 242523 251695 242529 251755
rect 242474 251683 242529 251695
rect 242641 251755 242694 251767
rect 242641 251695 242647 251755
rect 242681 251695 242694 251755
rect 242641 251683 242694 251695
rect 242474 251680 242508 251683
rect 242263 251645 242355 251651
rect 242263 251611 242275 251645
rect 242343 251611 242355 251645
rect 242263 251605 242355 251611
rect 242539 251645 242631 251651
rect 242539 251611 242551 251645
rect 242619 251611 242631 251645
rect 242539 251605 242631 251611
rect 242664 251518 242694 251683
rect 242752 251767 242782 251778
rect 242946 251767 242980 251942
rect 242752 251755 242805 251767
rect 242752 251695 242765 251755
rect 242799 251695 242805 251755
rect 242752 251683 242805 251695
rect 242917 251755 242980 251767
rect 242917 251695 242923 251755
rect 242957 251695 242980 251755
rect 242917 251683 242980 251695
rect 242752 251518 242782 251683
rect 242946 251678 242980 251683
rect 243024 251767 243058 251942
rect 243091 251839 243183 251845
rect 243091 251805 243103 251839
rect 243171 251805 243183 251839
rect 243091 251799 243183 251805
rect 243367 251839 243459 251845
rect 243367 251805 243379 251839
rect 243447 251805 243459 251839
rect 243367 251799 243459 251805
rect 243216 251767 243246 251782
rect 243024 251755 243081 251767
rect 243024 251695 243041 251755
rect 243075 251695 243081 251755
rect 243024 251683 243081 251695
rect 243193 251755 243246 251767
rect 243193 251695 243199 251755
rect 243233 251695 243246 251755
rect 243193 251683 243246 251695
rect 243024 251680 243058 251683
rect 242815 251645 242907 251651
rect 242815 251611 242827 251645
rect 242895 251611 242907 251645
rect 242815 251605 242907 251611
rect 243091 251645 243183 251651
rect 243091 251611 243103 251645
rect 243171 251611 243183 251645
rect 243091 251605 243183 251611
rect 243216 251518 243246 251683
rect 243304 251767 243334 251782
rect 243502 251767 243536 251942
rect 243304 251755 243357 251767
rect 243304 251695 243317 251755
rect 243351 251695 243357 251755
rect 243304 251683 243357 251695
rect 243469 251755 243536 251767
rect 243469 251695 243475 251755
rect 243509 251695 243536 251755
rect 243469 251683 243536 251695
rect 243304 251518 243334 251683
rect 243502 251670 243536 251683
rect 243576 251767 243610 251942
rect 243643 251839 243735 251845
rect 243643 251805 243655 251839
rect 243723 251805 243735 251839
rect 243643 251799 243735 251805
rect 243919 251839 244011 251845
rect 243919 251805 243931 251839
rect 243999 251805 244011 251839
rect 243919 251799 244011 251805
rect 243766 251767 243796 251784
rect 243576 251755 243633 251767
rect 243576 251695 243593 251755
rect 243627 251695 243633 251755
rect 243576 251683 243633 251695
rect 243745 251755 243796 251767
rect 243745 251695 243751 251755
rect 243785 251695 243796 251755
rect 243745 251683 243796 251695
rect 243576 251674 243610 251683
rect 243367 251645 243459 251651
rect 243367 251611 243379 251645
rect 243447 251611 243459 251645
rect 243367 251605 243459 251611
rect 243643 251645 243735 251651
rect 243643 251611 243655 251645
rect 243723 251611 243735 251645
rect 243643 251605 243735 251611
rect 243766 251518 243796 251683
rect 243854 251767 243884 251782
rect 244046 251767 244080 251942
rect 243854 251755 243909 251767
rect 243854 251695 243869 251755
rect 243903 251695 243909 251755
rect 243854 251683 243909 251695
rect 244021 251755 244080 251767
rect 244021 251695 244027 251755
rect 244061 251695 244080 251755
rect 244021 251683 244080 251695
rect 243854 251518 243884 251683
rect 244046 251670 244080 251683
rect 244126 251767 244160 251942
rect 244195 251839 244287 251845
rect 244195 251805 244207 251839
rect 244275 251805 244287 251839
rect 244195 251799 244287 251805
rect 244471 251839 244563 251845
rect 244471 251805 244483 251839
rect 244551 251805 244563 251839
rect 244471 251799 244563 251805
rect 244318 251767 244348 251782
rect 244126 251755 244185 251767
rect 244126 251695 244145 251755
rect 244179 251695 244185 251755
rect 244126 251683 244185 251695
rect 244297 251755 244348 251767
rect 244297 251695 244303 251755
rect 244337 251695 244348 251755
rect 244297 251683 244348 251695
rect 244126 251668 244160 251683
rect 243919 251645 244011 251651
rect 243919 251611 243931 251645
rect 243999 251611 244011 251645
rect 243919 251605 244011 251611
rect 244195 251645 244287 251651
rect 244195 251611 244207 251645
rect 244275 251611 244287 251645
rect 244195 251605 244287 251611
rect 244318 251518 244348 251683
rect 244406 251767 244436 251784
rect 244602 251767 244636 251942
rect 244406 251755 244461 251767
rect 244406 251695 244421 251755
rect 244455 251695 244461 251755
rect 244406 251683 244461 251695
rect 244573 251755 244636 251767
rect 244573 251695 244579 251755
rect 244613 251695 244636 251755
rect 244573 251683 244636 251695
rect 244406 251518 244436 251683
rect 244602 251670 244636 251683
rect 244676 251767 244710 251942
rect 244747 251839 244839 251845
rect 244747 251805 244759 251839
rect 244827 251805 244839 251839
rect 244747 251799 244839 251805
rect 245023 251839 245115 251845
rect 245023 251805 245035 251839
rect 245103 251805 245115 251839
rect 245023 251799 245115 251805
rect 244870 251767 244900 251782
rect 244676 251755 244737 251767
rect 244676 251695 244697 251755
rect 244731 251695 244737 251755
rect 244676 251683 244737 251695
rect 244849 251755 244900 251767
rect 244849 251695 244855 251755
rect 244889 251695 244900 251755
rect 244849 251683 244900 251695
rect 244676 251668 244710 251683
rect 244471 251645 244563 251651
rect 244471 251611 244483 251645
rect 244551 251611 244563 251645
rect 244471 251605 244563 251611
rect 244747 251645 244839 251651
rect 244747 251611 244759 251645
rect 244827 251611 244839 251645
rect 244747 251605 244839 251611
rect 244870 251518 244900 251683
rect 244960 251767 244990 251784
rect 245152 251767 245186 251942
rect 244960 251755 245013 251767
rect 244960 251695 244973 251755
rect 245007 251695 245013 251755
rect 244960 251683 245013 251695
rect 245125 251755 245186 251767
rect 245125 251695 245131 251755
rect 245165 251695 245186 251755
rect 245125 251683 245186 251695
rect 244960 251518 244990 251683
rect 245152 251672 245186 251683
rect 245228 251767 245262 251942
rect 245299 251839 245391 251845
rect 245299 251805 245311 251839
rect 245379 251805 245391 251839
rect 245299 251799 245391 251805
rect 245575 251839 245667 251845
rect 245575 251805 245587 251839
rect 245655 251805 245667 251839
rect 245575 251799 245667 251805
rect 245422 251767 245452 251782
rect 245228 251755 245289 251767
rect 245228 251695 245249 251755
rect 245283 251695 245289 251755
rect 245228 251683 245289 251695
rect 245401 251755 245452 251767
rect 245401 251695 245407 251755
rect 245441 251695 245452 251755
rect 245401 251683 245452 251695
rect 245228 251672 245262 251683
rect 245023 251645 245115 251651
rect 245023 251611 245035 251645
rect 245103 251611 245115 251645
rect 245023 251605 245115 251611
rect 245299 251645 245391 251651
rect 245299 251611 245311 251645
rect 245379 251611 245391 251645
rect 245299 251605 245391 251611
rect 245422 251518 245452 251683
rect 245512 251767 245542 251784
rect 245702 251767 245736 251942
rect 245512 251755 245565 251767
rect 245512 251695 245525 251755
rect 245559 251695 245565 251755
rect 245512 251683 245565 251695
rect 245677 251755 245736 251767
rect 245677 251695 245683 251755
rect 245717 251695 245736 251755
rect 245677 251683 245736 251695
rect 245512 251518 245542 251683
rect 245702 251676 245736 251683
rect 245784 251767 245818 251942
rect 245851 251839 245943 251845
rect 245851 251805 245863 251839
rect 245931 251805 245943 251839
rect 245851 251799 245943 251805
rect 246127 251839 246219 251845
rect 246127 251805 246139 251839
rect 246207 251805 246219 251839
rect 246127 251799 246219 251805
rect 245976 251767 246006 251788
rect 245784 251755 245841 251767
rect 245784 251695 245801 251755
rect 245835 251695 245841 251755
rect 245784 251683 245841 251695
rect 245953 251755 246006 251767
rect 245953 251695 245959 251755
rect 245993 251695 246006 251755
rect 245953 251683 246006 251695
rect 245784 251674 245818 251683
rect 245575 251645 245667 251651
rect 245575 251611 245587 251645
rect 245655 251611 245667 251645
rect 245575 251605 245667 251611
rect 245851 251645 245943 251651
rect 245851 251611 245863 251645
rect 245931 251611 245943 251645
rect 245851 251605 245943 251611
rect 245976 251518 246006 251683
rect 246066 251767 246096 251790
rect 246254 251767 246288 251942
rect 246066 251755 246117 251767
rect 246066 251695 246077 251755
rect 246111 251695 246117 251755
rect 246066 251683 246117 251695
rect 246229 251755 246288 251767
rect 246229 251695 246235 251755
rect 246269 251695 246288 251755
rect 246229 251683 246288 251695
rect 246066 251518 246096 251683
rect 246254 251680 246288 251683
rect 246332 251767 246366 251942
rect 246403 251839 246495 251845
rect 246403 251805 246415 251839
rect 246483 251805 246495 251839
rect 246403 251799 246495 251805
rect 246679 251839 246771 251845
rect 246679 251805 246691 251839
rect 246759 251805 246771 251839
rect 246679 251799 246771 251805
rect 246530 251767 246560 251790
rect 246332 251755 246393 251767
rect 246332 251695 246353 251755
rect 246387 251695 246393 251755
rect 246332 251683 246393 251695
rect 246505 251755 246560 251767
rect 246505 251695 246511 251755
rect 246545 251695 246560 251755
rect 246505 251683 246560 251695
rect 246332 251682 246366 251683
rect 246127 251645 246219 251651
rect 246127 251611 246139 251645
rect 246207 251611 246219 251645
rect 246127 251605 246219 251611
rect 246403 251645 246495 251651
rect 246403 251611 246415 251645
rect 246483 251611 246495 251645
rect 246403 251605 246495 251611
rect 246530 251518 246560 251683
rect 246616 251767 246646 251794
rect 246804 251767 246838 251942
rect 246616 251755 246669 251767
rect 246616 251695 246629 251755
rect 246663 251695 246669 251755
rect 246616 251683 246669 251695
rect 246781 251755 246838 251767
rect 246781 251695 246787 251755
rect 246821 251695 246838 251755
rect 246781 251683 246838 251695
rect 246616 251518 246646 251683
rect 246804 251678 246838 251683
rect 246888 251767 246922 251942
rect 246955 251839 247047 251845
rect 246955 251805 246967 251839
rect 247035 251805 247047 251839
rect 246955 251799 247047 251805
rect 247231 251839 247323 251845
rect 247231 251805 247243 251839
rect 247311 251805 247323 251839
rect 247231 251799 247323 251805
rect 247076 251767 247106 251780
rect 246888 251755 246945 251767
rect 246888 251695 246905 251755
rect 246939 251695 246945 251755
rect 246888 251683 246945 251695
rect 247057 251755 247106 251767
rect 247057 251695 247063 251755
rect 247097 251695 247106 251755
rect 247057 251683 247106 251695
rect 246888 251676 246922 251683
rect 246679 251645 246771 251651
rect 246679 251611 246691 251645
rect 246759 251611 246771 251645
rect 246679 251605 246771 251611
rect 246955 251645 247047 251651
rect 246955 251611 246967 251645
rect 247035 251611 247047 251645
rect 246955 251605 247047 251611
rect 247076 251518 247106 251683
rect 247168 251767 247198 251778
rect 247356 251767 247390 251942
rect 247168 251755 247221 251767
rect 247168 251695 247181 251755
rect 247215 251695 247221 251755
rect 247168 251683 247221 251695
rect 247333 251755 247390 251767
rect 247333 251695 247339 251755
rect 247373 251695 247390 251755
rect 247333 251683 247390 251695
rect 247168 251518 247198 251683
rect 247356 251678 247390 251683
rect 247440 251767 247474 251942
rect 247507 251839 247599 251845
rect 247507 251805 247519 251839
rect 247587 251805 247599 251839
rect 247507 251799 247599 251805
rect 247783 251839 247875 251845
rect 247783 251805 247795 251839
rect 247863 251805 247875 251839
rect 247783 251799 247875 251805
rect 247632 251767 247662 251780
rect 247440 251755 247497 251767
rect 247440 251695 247457 251755
rect 247491 251695 247497 251755
rect 247440 251683 247497 251695
rect 247609 251755 247662 251767
rect 247609 251695 247615 251755
rect 247649 251695 247662 251755
rect 247609 251683 247662 251695
rect 247440 251680 247474 251683
rect 247231 251645 247323 251651
rect 247231 251611 247243 251645
rect 247311 251611 247323 251645
rect 247231 251605 247323 251611
rect 247507 251645 247599 251651
rect 247507 251611 247519 251645
rect 247587 251611 247599 251645
rect 247507 251605 247599 251611
rect 247632 251518 247662 251683
rect 247716 251767 247746 251780
rect 247910 251767 247944 251942
rect 247716 251755 247773 251767
rect 247716 251695 247733 251755
rect 247767 251695 247773 251755
rect 247716 251683 247773 251695
rect 247885 251755 247944 251767
rect 247885 251695 247891 251755
rect 247925 251695 247944 251755
rect 247885 251684 247944 251695
rect 247988 251767 248022 251942
rect 248059 251839 248151 251845
rect 248059 251805 248071 251839
rect 248139 251805 248151 251839
rect 248059 251799 248151 251805
rect 248182 251767 248212 251780
rect 247988 251755 248049 251767
rect 247988 251695 248009 251755
rect 248043 251695 248049 251755
rect 247885 251683 247931 251684
rect 247988 251683 248049 251695
rect 248161 251755 248212 251767
rect 248161 251695 248167 251755
rect 248201 251695 248212 251755
rect 248161 251683 248212 251695
rect 248302 251690 248336 251942
rect 247716 251518 247746 251683
rect 247988 251682 248022 251683
rect 247783 251645 247875 251651
rect 247783 251611 247795 251645
rect 247863 251611 247875 251645
rect 247783 251605 247875 251611
rect 248059 251645 248151 251651
rect 248059 251611 248071 251645
rect 248139 251611 248151 251645
rect 248059 251605 248151 251611
rect 248182 251518 248212 251683
rect 234045 251476 248214 251518
rect 248172 251474 248214 251476
rect 151792 251414 151992 251434
rect 238224 251370 238364 251382
rect 234266 251294 234350 251326
rect 234266 251252 234282 251294
rect 234336 251252 234350 251294
rect 147163 251184 150656 251230
rect 150154 251182 150186 251184
rect 59015 251172 60273 251174
rect 59017 251142 60273 251172
rect 234266 251164 234350 251252
rect 59017 251141 59585 251142
rect 59017 251138 59051 251141
rect 59293 251140 59585 251141
rect 148662 251130 148784 251140
rect 148662 251086 148690 251130
rect 148762 251086 148784 251130
rect 234266 251108 234274 251164
rect 234342 251108 234350 251164
rect 234266 251100 234350 251108
rect 238224 251314 238264 251370
rect 238342 251314 238364 251370
rect 58873 251044 59073 251066
rect 58812 250882 59076 251044
rect 59395 250996 59573 251026
rect 52872 250618 59076 250882
rect 59388 250990 59573 250996
rect 59388 250930 59439 250990
rect 59533 250930 59573 250990
rect 59388 250760 59573 250930
rect 148662 250904 148784 251086
rect 149124 251066 149214 251082
rect 149124 251002 149136 251066
rect 149208 251002 149214 251066
rect 148628 250896 148828 250904
rect 52872 249146 53136 250618
rect 59388 250340 59564 250760
rect 147552 250704 148828 250896
rect 147552 250678 148826 250704
rect 141996 250632 148826 250678
rect 141996 250414 147816 250632
rect 57078 249740 61758 250340
rect 52310 240230 53762 249146
rect 57078 248820 58038 249740
rect 57078 248220 57238 248820
rect 57838 248220 58038 248820
rect 57078 248060 58038 248220
rect 60798 248820 61758 249740
rect 141996 248942 142260 250414
rect 149124 250136 149214 251002
rect 238224 250700 238364 251314
rect 249168 251218 249968 251942
rect 249168 250972 249238 251218
rect 249378 250972 249968 251218
rect 249168 250886 249968 250972
rect 320433 250873 321381 251842
rect 411258 251469 412348 252005
rect 428318 251723 429188 251755
rect 413461 251657 429188 251723
rect 413341 251553 413433 251559
rect 413341 251519 413353 251553
rect 413421 251519 413433 251553
rect 413341 251513 413433 251519
rect 413466 251481 413506 251657
rect 413285 251469 413331 251481
rect 411258 251411 413291 251469
rect 337608 251127 339092 251157
rect 322818 251061 339092 251127
rect 322698 250957 322790 250963
rect 322698 250923 322710 250957
rect 322778 250923 322790 250957
rect 322698 250917 322790 250923
rect 322823 250885 322863 251061
rect 322642 250873 322688 250885
rect 320433 250815 322648 250873
rect 320433 250798 321381 250815
rect 233248 250500 238410 250700
rect 322484 250637 322526 250815
rect 322642 250813 322648 250815
rect 322682 250813 322688 250873
rect 322642 250801 322688 250813
rect 322800 250873 322863 250885
rect 322800 250813 322806 250873
rect 322840 250813 322863 250873
rect 322800 250801 322863 250813
rect 322823 250795 322863 250801
rect 322905 250885 322945 251061
rect 322974 250957 323066 250963
rect 322974 250923 322986 250957
rect 323054 250923 323066 250957
rect 322974 250917 323066 250923
rect 323250 250957 323342 250963
rect 323250 250923 323262 250957
rect 323330 250923 323342 250957
rect 323250 250917 323342 250923
rect 323099 250885 323129 250893
rect 322905 250873 322964 250885
rect 322905 250813 322924 250873
rect 322958 250813 322964 250873
rect 322905 250801 322964 250813
rect 323076 250873 323129 250885
rect 323076 250813 323082 250873
rect 323116 250813 323129 250873
rect 323076 250801 323129 250813
rect 322905 250797 322945 250801
rect 322698 250763 322790 250769
rect 322698 250729 322710 250763
rect 322778 250729 322790 250763
rect 322698 250723 322790 250729
rect 322974 250763 323066 250769
rect 322974 250729 322986 250763
rect 323054 250729 323066 250763
rect 322974 250723 323066 250729
rect 323099 250637 323129 250801
rect 323185 250885 323215 250893
rect 323381 250885 323421 251061
rect 323185 250873 323240 250885
rect 323185 250813 323200 250873
rect 323234 250813 323240 250873
rect 323185 250801 323240 250813
rect 323352 250873 323421 250885
rect 323352 250813 323358 250873
rect 323392 250813 323421 250873
rect 323352 250801 323421 250813
rect 323185 250637 323215 250801
rect 323381 250797 323421 250801
rect 323449 250885 323489 251061
rect 323526 250957 323618 250963
rect 323526 250923 323538 250957
rect 323606 250923 323618 250957
rect 323526 250917 323618 250923
rect 323802 250957 323894 250963
rect 323802 250923 323814 250957
rect 323882 250923 323894 250957
rect 323802 250917 323894 250923
rect 323653 250885 323683 250893
rect 323449 250873 323516 250885
rect 323449 250813 323476 250873
rect 323510 250813 323516 250873
rect 323449 250801 323516 250813
rect 323628 250873 323683 250885
rect 323628 250813 323634 250873
rect 323668 250813 323683 250873
rect 323628 250801 323683 250813
rect 323449 250797 323489 250801
rect 323250 250763 323342 250769
rect 323250 250729 323262 250763
rect 323330 250729 323342 250763
rect 323250 250723 323342 250729
rect 323526 250763 323618 250769
rect 323526 250729 323538 250763
rect 323606 250729 323618 250763
rect 323526 250723 323618 250729
rect 323653 250637 323683 250801
rect 323739 250885 323769 250893
rect 323929 250885 323969 251061
rect 323739 250873 323792 250885
rect 323739 250813 323752 250873
rect 323786 250813 323792 250873
rect 323739 250801 323792 250813
rect 323904 250873 323969 250885
rect 323904 250813 323910 250873
rect 323944 250813 323969 250873
rect 323904 250801 323969 250813
rect 323739 250637 323769 250801
rect 323929 250793 323969 250801
rect 324001 250885 324041 251061
rect 324078 250957 324170 250963
rect 324078 250923 324090 250957
rect 324158 250923 324170 250957
rect 324078 250917 324170 250923
rect 324354 250957 324446 250963
rect 324354 250923 324366 250957
rect 324434 250923 324446 250957
rect 324354 250917 324446 250923
rect 324201 250885 324231 250893
rect 324001 250873 324068 250885
rect 324001 250813 324028 250873
rect 324062 250813 324068 250873
rect 324001 250801 324068 250813
rect 324180 250873 324231 250885
rect 324180 250813 324186 250873
rect 324220 250813 324231 250873
rect 324180 250801 324231 250813
rect 324001 250797 324041 250801
rect 323802 250763 323894 250769
rect 323802 250729 323814 250763
rect 323882 250729 323894 250763
rect 323802 250723 323894 250729
rect 324078 250763 324170 250769
rect 324078 250729 324090 250763
rect 324158 250729 324170 250763
rect 324078 250723 324170 250729
rect 324201 250637 324231 250801
rect 324293 250885 324323 250891
rect 324481 250885 324521 251061
rect 324293 250873 324344 250885
rect 324293 250813 324304 250873
rect 324338 250813 324344 250873
rect 324293 250801 324344 250813
rect 324456 250873 324521 250885
rect 324456 250813 324462 250873
rect 324496 250813 324521 250873
rect 324456 250801 324521 250813
rect 324561 250885 324601 251061
rect 324630 250957 324722 250963
rect 324630 250923 324642 250957
rect 324710 250923 324722 250957
rect 324630 250917 324722 250923
rect 324906 250957 324998 250963
rect 324906 250923 324918 250957
rect 324986 250923 324998 250957
rect 324906 250917 324998 250923
rect 324751 250885 324781 250891
rect 324561 250873 324620 250885
rect 324561 250813 324580 250873
rect 324614 250813 324620 250873
rect 324561 250801 324620 250813
rect 324732 250873 324781 250885
rect 324732 250813 324738 250873
rect 324772 250813 324781 250873
rect 324732 250801 324781 250813
rect 324293 250637 324323 250801
rect 324354 250763 324446 250769
rect 324354 250729 324366 250763
rect 324434 250729 324446 250763
rect 324354 250723 324446 250729
rect 324630 250763 324722 250769
rect 324630 250729 324642 250763
rect 324710 250729 324722 250763
rect 324630 250723 324722 250729
rect 324751 250637 324781 250801
rect 324843 250885 324873 250889
rect 325035 250885 325075 251061
rect 324843 250873 324896 250885
rect 324843 250813 324856 250873
rect 324890 250813 324896 250873
rect 324843 250801 324896 250813
rect 325008 250873 325075 250885
rect 325008 250813 325014 250873
rect 325048 250813 325075 250873
rect 325008 250801 325075 250813
rect 324843 250637 324873 250801
rect 325035 250797 325075 250801
rect 325109 250885 325149 251061
rect 325182 250957 325274 250963
rect 325182 250923 325194 250957
rect 325262 250923 325274 250957
rect 325182 250917 325274 250923
rect 325458 250957 325550 250963
rect 325458 250923 325470 250957
rect 325538 250923 325550 250957
rect 325458 250917 325550 250923
rect 325307 250885 325337 250889
rect 325109 250873 325172 250885
rect 325109 250813 325132 250873
rect 325166 250813 325172 250873
rect 325109 250801 325172 250813
rect 325284 250873 325337 250885
rect 325284 250813 325290 250873
rect 325324 250813 325337 250873
rect 325284 250801 325337 250813
rect 325109 250799 325149 250801
rect 324906 250763 324998 250769
rect 324906 250729 324918 250763
rect 324986 250729 324998 250763
rect 324906 250723 324998 250729
rect 325182 250763 325274 250769
rect 325182 250729 325194 250763
rect 325262 250729 325274 250763
rect 325182 250723 325274 250729
rect 325307 250637 325337 250801
rect 325395 250885 325425 250887
rect 325587 250885 325627 251061
rect 325395 250873 325448 250885
rect 325395 250813 325408 250873
rect 325442 250813 325448 250873
rect 325395 250801 325448 250813
rect 325560 250873 325627 250885
rect 325560 250813 325566 250873
rect 325600 250813 325627 250873
rect 325560 250801 325627 250813
rect 325395 250637 325425 250801
rect 325587 250795 325627 250801
rect 325657 250885 325697 251061
rect 325734 250957 325826 250963
rect 325734 250923 325746 250957
rect 325814 250923 325826 250957
rect 325734 250917 325826 250923
rect 326010 250957 326102 250963
rect 326010 250923 326022 250957
rect 326090 250923 326102 250957
rect 326010 250917 326102 250923
rect 325857 250885 325887 250887
rect 325657 250873 325724 250885
rect 325657 250813 325684 250873
rect 325718 250813 325724 250873
rect 325657 250801 325724 250813
rect 325836 250873 325887 250885
rect 325836 250813 325842 250873
rect 325876 250813 325887 250873
rect 325836 250801 325887 250813
rect 325657 250799 325697 250801
rect 325458 250763 325550 250769
rect 325734 250767 325826 250769
rect 325458 250729 325470 250763
rect 325538 250729 325550 250763
rect 325731 250763 325826 250767
rect 325731 250734 325746 250763
rect 325458 250723 325550 250729
rect 325734 250729 325746 250734
rect 325814 250729 325826 250763
rect 325734 250723 325826 250729
rect 325857 250637 325887 250801
rect 325945 250885 325975 250887
rect 326135 250885 326175 251061
rect 325945 250873 326000 250885
rect 325945 250813 325960 250873
rect 325994 250813 326000 250873
rect 325945 250801 326000 250813
rect 326112 250873 326175 250885
rect 326112 250813 326118 250873
rect 326152 250813 326175 250873
rect 326112 250801 326175 250813
rect 325945 250637 325975 250801
rect 326135 250795 326175 250801
rect 326213 250885 326253 251061
rect 326286 250957 326378 250963
rect 326286 250923 326298 250957
rect 326366 250923 326378 250957
rect 326286 250917 326378 250923
rect 326562 250957 326654 250963
rect 326562 250923 326574 250957
rect 326642 250923 326654 250957
rect 326562 250917 326654 250923
rect 326409 250885 326439 250889
rect 326213 250873 326276 250885
rect 326213 250813 326236 250873
rect 326270 250813 326276 250873
rect 326213 250801 326276 250813
rect 326388 250873 326439 250885
rect 326388 250813 326394 250873
rect 326428 250813 326439 250873
rect 326388 250801 326439 250813
rect 326213 250799 326253 250801
rect 326010 250763 326102 250769
rect 326010 250729 326022 250763
rect 326090 250729 326102 250763
rect 326010 250723 326102 250729
rect 326286 250763 326378 250769
rect 326286 250729 326298 250763
rect 326366 250729 326378 250763
rect 326286 250723 326378 250729
rect 326409 250637 326439 250801
rect 326497 250885 326527 250889
rect 326689 250885 326729 251061
rect 326497 250873 326552 250885
rect 326497 250813 326512 250873
rect 326546 250813 326552 250873
rect 326497 250801 326552 250813
rect 326664 250873 326729 250885
rect 326664 250813 326670 250873
rect 326704 250813 326729 250873
rect 326664 250801 326729 250813
rect 326497 250637 326527 250801
rect 326689 250787 326729 250801
rect 326767 250885 326807 251061
rect 326838 250957 326930 250963
rect 326838 250923 326850 250957
rect 326918 250923 326930 250957
rect 326838 250917 326930 250923
rect 327114 250957 327206 250963
rect 327114 250923 327126 250957
rect 327194 250923 327206 250957
rect 327114 250917 327206 250923
rect 326961 250885 326991 250889
rect 326767 250873 326828 250885
rect 326767 250813 326788 250873
rect 326822 250813 326828 250873
rect 326767 250801 326828 250813
rect 326940 250873 326991 250885
rect 326940 250813 326946 250873
rect 326980 250813 326991 250873
rect 326940 250801 326991 250813
rect 326767 250795 326807 250801
rect 326562 250763 326654 250769
rect 326562 250729 326574 250763
rect 326642 250729 326654 250763
rect 326562 250723 326654 250729
rect 326838 250763 326930 250769
rect 326838 250729 326850 250763
rect 326918 250729 326930 250763
rect 326838 250723 326930 250729
rect 326961 250637 326991 250801
rect 327053 250885 327083 250889
rect 327245 250885 327285 251061
rect 327053 250873 327104 250885
rect 327053 250813 327064 250873
rect 327098 250813 327104 250873
rect 327053 250801 327104 250813
rect 327216 250873 327285 250885
rect 327216 250813 327222 250873
rect 327256 250813 327285 250873
rect 327216 250801 327285 250813
rect 327319 250885 327359 251061
rect 327390 250957 327482 250963
rect 327390 250923 327402 250957
rect 327470 250923 327482 250957
rect 327390 250917 327482 250923
rect 327666 250957 327758 250963
rect 327666 250923 327678 250957
rect 327746 250923 327758 250957
rect 327666 250917 327758 250923
rect 327515 250885 327545 250899
rect 327319 250873 327380 250885
rect 327319 250813 327340 250873
rect 327374 250813 327380 250873
rect 327319 250801 327380 250813
rect 327492 250873 327545 250885
rect 327492 250813 327498 250873
rect 327532 250813 327545 250873
rect 327492 250801 327545 250813
rect 327053 250637 327083 250801
rect 327245 250797 327285 250801
rect 327114 250763 327206 250769
rect 327114 250729 327126 250763
rect 327194 250729 327206 250763
rect 327114 250723 327206 250729
rect 327390 250763 327482 250769
rect 327390 250729 327402 250763
rect 327470 250729 327482 250763
rect 327390 250723 327482 250729
rect 327515 250637 327545 250801
rect 327601 250885 327631 250897
rect 327789 250885 327823 251061
rect 327601 250873 327656 250885
rect 327601 250813 327616 250873
rect 327650 250813 327656 250873
rect 327601 250801 327656 250813
rect 327768 250873 327823 250885
rect 327768 250813 327774 250873
rect 327808 250813 327823 250873
rect 327768 250801 327823 250813
rect 327601 250637 327631 250801
rect 327789 250797 327823 250801
rect 327879 250885 327913 251061
rect 327942 250957 328034 250963
rect 327942 250923 327954 250957
rect 328022 250923 328034 250957
rect 327942 250917 328034 250923
rect 328218 250957 328310 250963
rect 328218 250923 328230 250957
rect 328298 250923 328310 250957
rect 328218 250917 328310 250923
rect 328069 250885 328099 250895
rect 327879 250873 327932 250885
rect 327879 250813 327892 250873
rect 327926 250813 327932 250873
rect 327879 250801 327932 250813
rect 328044 250873 328099 250885
rect 328044 250813 328050 250873
rect 328084 250813 328099 250873
rect 328044 250801 328099 250813
rect 327879 250797 327913 250801
rect 327666 250763 327758 250769
rect 327666 250729 327678 250763
rect 327746 250729 327758 250763
rect 327666 250723 327758 250729
rect 327942 250763 328034 250769
rect 327942 250729 327954 250763
rect 328022 250729 328034 250763
rect 327942 250723 328034 250729
rect 328069 250637 328099 250801
rect 328155 250885 328185 250895
rect 328345 250885 328379 251061
rect 328155 250873 328208 250885
rect 328155 250813 328168 250873
rect 328202 250813 328208 250873
rect 328155 250801 328208 250813
rect 328320 250873 328379 250885
rect 328320 250813 328326 250873
rect 328360 250813 328379 250873
rect 328320 250801 328379 250813
rect 328429 250885 328463 251061
rect 328494 250957 328586 250963
rect 328494 250923 328506 250957
rect 328574 250923 328586 250957
rect 328494 250917 328586 250923
rect 328621 250885 328655 250899
rect 328429 250873 328484 250885
rect 328429 250813 328444 250873
rect 328478 250813 328484 250873
rect 328429 250801 328484 250813
rect 328596 250873 328655 250885
rect 328596 250813 328602 250873
rect 328636 250813 328655 250873
rect 328596 250801 328655 250813
rect 328155 250637 328185 250801
rect 328345 250797 328379 250801
rect 328218 250763 328310 250769
rect 328218 250729 328230 250763
rect 328298 250729 328310 250763
rect 328218 250723 328310 250729
rect 328494 250763 328586 250769
rect 328494 250729 328506 250763
rect 328574 250729 328586 250763
rect 328494 250723 328586 250729
rect 328621 250637 328655 250801
rect 328703 250885 328737 251061
rect 328770 250957 328862 250963
rect 328770 250923 328782 250957
rect 328850 250923 328862 250957
rect 328770 250917 328862 250923
rect 329046 250957 329138 250963
rect 329046 250923 329058 250957
rect 329126 250923 329138 250957
rect 329046 250917 329138 250923
rect 328895 250885 328925 250897
rect 328703 250873 328760 250885
rect 328703 250813 328720 250873
rect 328754 250813 328760 250873
rect 328703 250801 328760 250813
rect 328872 250873 328925 250885
rect 328872 250813 328878 250873
rect 328912 250813 328925 250873
rect 328872 250801 328925 250813
rect 328703 250799 328737 250801
rect 328770 250763 328862 250769
rect 328770 250729 328782 250763
rect 328850 250729 328862 250763
rect 328770 250723 328862 250729
rect 328895 250637 328925 250801
rect 328983 250885 329013 250899
rect 329173 250885 329207 251061
rect 328983 250873 329036 250885
rect 328983 250813 328996 250873
rect 329030 250813 329036 250873
rect 328983 250801 329036 250813
rect 329148 250873 329207 250885
rect 329148 250813 329154 250873
rect 329188 250813 329207 250873
rect 329148 250801 329207 250813
rect 329259 250885 329293 251061
rect 329331 250999 329546 251009
rect 329331 250963 329461 250999
rect 329322 250957 329461 250963
rect 329322 250923 329334 250957
rect 329402 250939 329461 250957
rect 329521 250939 329546 250999
rect 329402 250929 329546 250939
rect 329598 250957 329690 250963
rect 329402 250923 329414 250929
rect 329322 250917 329414 250923
rect 329598 250923 329610 250957
rect 329678 250923 329690 250957
rect 329598 250917 329690 250923
rect 329443 250885 329473 250899
rect 329259 250873 329312 250885
rect 329259 250813 329272 250873
rect 329306 250813 329312 250873
rect 329259 250801 329312 250813
rect 329424 250873 329473 250885
rect 329424 250813 329430 250873
rect 329464 250813 329473 250873
rect 329424 250801 329473 250813
rect 328983 250637 329013 250801
rect 329259 250795 329293 250801
rect 329046 250763 329138 250769
rect 329046 250729 329058 250763
rect 329126 250729 329138 250763
rect 329322 250763 329414 250769
rect 329322 250744 329334 250763
rect 329046 250723 329138 250729
rect 329186 250739 329334 250744
rect 329186 250684 329196 250739
rect 329261 250729 329334 250739
rect 329402 250729 329414 250763
rect 329261 250723 329414 250729
rect 329261 250694 329401 250723
rect 329261 250684 329271 250694
rect 329186 250679 329271 250684
rect 329443 250637 329473 250801
rect 329535 250885 329565 250899
rect 329725 250885 329759 251061
rect 329535 250873 329588 250885
rect 329535 250813 329548 250873
rect 329582 250813 329588 250873
rect 329535 250801 329588 250813
rect 329700 250873 329759 250885
rect 329700 250813 329706 250873
rect 329740 250813 329759 250873
rect 329700 250803 329759 250813
rect 329811 250885 329845 251061
rect 329874 250957 329966 250963
rect 329874 250923 329886 250957
rect 329954 250923 329966 250957
rect 329874 250917 329966 250923
rect 330150 250957 330242 250963
rect 330150 250923 330162 250957
rect 330230 250923 330242 250957
rect 330150 250917 330242 250923
rect 329997 250885 330027 250899
rect 329811 250873 329864 250885
rect 329811 250813 329824 250873
rect 329858 250813 329864 250873
rect 329700 250801 329746 250803
rect 329811 250801 329864 250813
rect 329976 250873 330027 250885
rect 329976 250813 329982 250873
rect 330016 250813 330027 250873
rect 329976 250801 330027 250813
rect 329535 250637 329565 250801
rect 329811 250799 329845 250801
rect 329598 250763 329690 250769
rect 329598 250729 329610 250763
rect 329678 250729 329690 250763
rect 329598 250723 329690 250729
rect 329874 250763 329966 250769
rect 329874 250729 329886 250763
rect 329954 250729 329966 250763
rect 329874 250723 329966 250729
rect 329997 250637 330027 250801
rect 330089 250885 330119 250899
rect 330275 250885 330309 251061
rect 330089 250873 330140 250885
rect 330089 250813 330100 250873
rect 330134 250813 330140 250873
rect 330089 250801 330140 250813
rect 330252 250873 330309 250885
rect 330252 250813 330258 250873
rect 330292 250813 330309 250873
rect 330252 250801 330309 250813
rect 330089 250637 330119 250801
rect 330275 250799 330309 250801
rect 330363 250885 330397 251061
rect 330426 250957 330518 250963
rect 330426 250923 330438 250957
rect 330506 250923 330518 250957
rect 330426 250917 330518 250923
rect 330702 250957 330794 250963
rect 330702 250923 330714 250957
rect 330782 250923 330794 250957
rect 330702 250917 330794 250923
rect 330549 250885 330579 250899
rect 330363 250873 330416 250885
rect 330363 250813 330376 250873
rect 330410 250813 330416 250873
rect 330363 250801 330416 250813
rect 330528 250873 330579 250885
rect 330528 250813 330534 250873
rect 330568 250813 330579 250873
rect 330528 250801 330579 250813
rect 330363 250797 330397 250801
rect 330150 250763 330242 250769
rect 330150 250729 330162 250763
rect 330230 250729 330242 250763
rect 330150 250723 330242 250729
rect 330426 250763 330518 250769
rect 330426 250729 330438 250763
rect 330506 250729 330518 250763
rect 330426 250723 330518 250729
rect 330549 250637 330579 250801
rect 330635 250885 330665 250899
rect 330831 250885 330865 251061
rect 330635 250873 330692 250885
rect 330635 250813 330652 250873
rect 330686 250813 330692 250873
rect 330635 250801 330692 250813
rect 330804 250873 330865 250885
rect 330804 250813 330810 250873
rect 330844 250813 330865 250873
rect 330804 250801 330865 250813
rect 330635 250637 330665 250801
rect 330831 250793 330865 250801
rect 330913 250885 330947 251061
rect 330978 250957 331070 250963
rect 330978 250923 330990 250957
rect 331058 250923 331070 250957
rect 330978 250917 331070 250923
rect 331254 250957 331346 250963
rect 331254 250923 331266 250957
rect 331334 250923 331346 250957
rect 331254 250917 331346 250923
rect 331103 250885 331133 250899
rect 330913 250873 330968 250885
rect 330913 250813 330928 250873
rect 330962 250813 330968 250873
rect 330913 250801 330968 250813
rect 331080 250873 331133 250885
rect 331080 250813 331086 250873
rect 331120 250813 331133 250873
rect 331080 250801 331133 250813
rect 330913 250799 330947 250801
rect 330702 250763 330794 250769
rect 330702 250729 330714 250763
rect 330782 250729 330794 250763
rect 330702 250723 330794 250729
rect 330978 250763 331070 250769
rect 330978 250729 330990 250763
rect 331058 250729 331070 250763
rect 330978 250723 331070 250729
rect 331103 250637 331133 250801
rect 331191 250885 331221 250897
rect 331385 250885 331419 251061
rect 331191 250873 331244 250885
rect 331191 250813 331204 250873
rect 331238 250813 331244 250873
rect 331191 250801 331244 250813
rect 331356 250873 331419 250885
rect 331356 250813 331362 250873
rect 331396 250813 331419 250873
rect 331356 250801 331419 250813
rect 331191 250637 331221 250801
rect 331385 250797 331419 250801
rect 331463 250885 331497 251061
rect 331530 250957 331622 250963
rect 331530 250923 331542 250957
rect 331610 250923 331622 250957
rect 331530 250917 331622 250923
rect 331806 250957 331898 250963
rect 331806 250923 331818 250957
rect 331886 250923 331898 250957
rect 331806 250917 331898 250923
rect 331655 250885 331685 250901
rect 331463 250873 331520 250885
rect 331463 250813 331480 250873
rect 331514 250813 331520 250873
rect 331463 250801 331520 250813
rect 331632 250873 331685 250885
rect 331632 250813 331638 250873
rect 331672 250813 331685 250873
rect 331632 250801 331685 250813
rect 331463 250799 331497 250801
rect 331254 250763 331346 250769
rect 331254 250729 331266 250763
rect 331334 250729 331346 250763
rect 331254 250723 331346 250729
rect 331530 250763 331622 250769
rect 331530 250729 331542 250763
rect 331610 250729 331622 250763
rect 331530 250723 331622 250729
rect 331655 250637 331685 250801
rect 331743 250885 331773 250901
rect 331941 250885 331975 251061
rect 331743 250873 331796 250885
rect 331743 250813 331756 250873
rect 331790 250813 331796 250873
rect 331743 250801 331796 250813
rect 331908 250873 331975 250885
rect 331908 250813 331914 250873
rect 331948 250813 331975 250873
rect 331908 250801 331975 250813
rect 331743 250637 331773 250801
rect 331941 250789 331975 250801
rect 332015 250885 332049 251061
rect 332082 250957 332174 250963
rect 332082 250923 332094 250957
rect 332162 250923 332174 250957
rect 332082 250917 332174 250923
rect 332358 250957 332450 250963
rect 332358 250923 332370 250957
rect 332438 250923 332450 250957
rect 332358 250917 332450 250923
rect 332205 250885 332235 250903
rect 332015 250873 332072 250885
rect 332015 250813 332032 250873
rect 332066 250813 332072 250873
rect 332015 250801 332072 250813
rect 332184 250873 332235 250885
rect 332184 250813 332190 250873
rect 332224 250813 332235 250873
rect 332184 250801 332235 250813
rect 332015 250793 332049 250801
rect 331806 250763 331898 250769
rect 331806 250729 331818 250763
rect 331886 250729 331898 250763
rect 331806 250723 331898 250729
rect 332082 250763 332174 250769
rect 332082 250729 332094 250763
rect 332162 250729 332174 250763
rect 332082 250723 332174 250729
rect 332205 250637 332235 250801
rect 332293 250885 332323 250901
rect 332485 250885 332519 251061
rect 332293 250873 332348 250885
rect 332293 250813 332308 250873
rect 332342 250813 332348 250873
rect 332293 250801 332348 250813
rect 332460 250873 332519 250885
rect 332460 250813 332466 250873
rect 332500 250813 332519 250873
rect 332460 250801 332519 250813
rect 332293 250637 332323 250801
rect 332485 250789 332519 250801
rect 332565 250885 332599 251061
rect 332634 250957 332726 250963
rect 332634 250923 332646 250957
rect 332714 250923 332726 250957
rect 332634 250917 332726 250923
rect 332910 250957 333002 250963
rect 332910 250923 332922 250957
rect 332990 250923 333002 250957
rect 332910 250917 333002 250923
rect 332757 250885 332787 250901
rect 332565 250873 332624 250885
rect 332565 250813 332584 250873
rect 332618 250813 332624 250873
rect 332565 250801 332624 250813
rect 332736 250873 332787 250885
rect 332736 250813 332742 250873
rect 332776 250813 332787 250873
rect 332736 250801 332787 250813
rect 332565 250787 332599 250801
rect 332358 250763 332450 250769
rect 332358 250729 332370 250763
rect 332438 250729 332450 250763
rect 332358 250723 332450 250729
rect 332634 250763 332726 250769
rect 332634 250729 332646 250763
rect 332714 250729 332726 250763
rect 332634 250723 332726 250729
rect 332757 250637 332787 250801
rect 332845 250885 332875 250903
rect 333041 250885 333075 251061
rect 332845 250873 332900 250885
rect 332845 250813 332860 250873
rect 332894 250813 332900 250873
rect 332845 250801 332900 250813
rect 333012 250873 333075 250885
rect 333012 250813 333018 250873
rect 333052 250813 333075 250873
rect 333012 250801 333075 250813
rect 332845 250637 332875 250801
rect 333041 250789 333075 250801
rect 333115 250885 333149 251061
rect 333186 250957 333278 250963
rect 333186 250923 333198 250957
rect 333266 250923 333278 250957
rect 333186 250917 333278 250923
rect 333462 250957 333554 250963
rect 333462 250923 333474 250957
rect 333542 250923 333554 250957
rect 333462 250917 333554 250923
rect 333309 250885 333339 250901
rect 333115 250873 333176 250885
rect 333115 250813 333136 250873
rect 333170 250813 333176 250873
rect 333115 250801 333176 250813
rect 333288 250873 333339 250885
rect 333288 250813 333294 250873
rect 333328 250813 333339 250873
rect 333288 250801 333339 250813
rect 333115 250787 333149 250801
rect 332910 250763 333002 250769
rect 332910 250729 332922 250763
rect 332990 250729 333002 250763
rect 332910 250723 333002 250729
rect 333186 250763 333278 250769
rect 333186 250729 333198 250763
rect 333266 250729 333278 250763
rect 333186 250723 333278 250729
rect 333309 250637 333339 250801
rect 333399 250885 333429 250903
rect 333591 250885 333625 251061
rect 333399 250873 333452 250885
rect 333399 250813 333412 250873
rect 333446 250813 333452 250873
rect 333399 250801 333452 250813
rect 333564 250873 333625 250885
rect 333564 250813 333570 250873
rect 333604 250813 333625 250873
rect 333564 250801 333625 250813
rect 333399 250637 333429 250801
rect 333591 250791 333625 250801
rect 333667 250885 333701 251061
rect 333738 250957 333830 250963
rect 333738 250923 333750 250957
rect 333818 250923 333830 250957
rect 333738 250917 333830 250923
rect 334014 250957 334106 250963
rect 334014 250923 334026 250957
rect 334094 250923 334106 250957
rect 334014 250917 334106 250923
rect 333861 250885 333891 250901
rect 333667 250873 333728 250885
rect 333667 250813 333688 250873
rect 333722 250813 333728 250873
rect 333667 250801 333728 250813
rect 333840 250873 333891 250885
rect 333840 250813 333846 250873
rect 333880 250813 333891 250873
rect 333840 250801 333891 250813
rect 333667 250791 333701 250801
rect 333462 250763 333554 250769
rect 333462 250729 333474 250763
rect 333542 250729 333554 250763
rect 333462 250723 333554 250729
rect 333738 250763 333830 250769
rect 333738 250729 333750 250763
rect 333818 250729 333830 250763
rect 333738 250723 333830 250729
rect 333861 250637 333891 250801
rect 333951 250885 333981 250903
rect 334141 250885 334175 251061
rect 333951 250873 334004 250885
rect 333951 250813 333964 250873
rect 333998 250813 334004 250873
rect 333951 250801 334004 250813
rect 334116 250873 334175 250885
rect 334116 250813 334122 250873
rect 334156 250813 334175 250873
rect 334116 250801 334175 250813
rect 333951 250637 333981 250801
rect 334141 250795 334175 250801
rect 334223 250885 334257 251061
rect 334290 250957 334382 250963
rect 334290 250923 334302 250957
rect 334370 250923 334382 250957
rect 334290 250917 334382 250923
rect 334566 250957 334658 250963
rect 334566 250923 334578 250957
rect 334646 250923 334658 250957
rect 334566 250917 334658 250923
rect 334415 250885 334445 250907
rect 334223 250873 334280 250885
rect 334223 250813 334240 250873
rect 334274 250813 334280 250873
rect 334223 250801 334280 250813
rect 334392 250873 334445 250885
rect 334392 250813 334398 250873
rect 334432 250813 334445 250873
rect 334392 250801 334445 250813
rect 334223 250793 334257 250801
rect 334014 250763 334106 250769
rect 334014 250729 334026 250763
rect 334094 250729 334106 250763
rect 334014 250723 334106 250729
rect 334290 250763 334382 250769
rect 334290 250729 334302 250763
rect 334370 250729 334382 250763
rect 334290 250723 334382 250729
rect 334415 250637 334445 250801
rect 334505 250885 334535 250909
rect 334693 250885 334727 251061
rect 334505 250873 334556 250885
rect 334505 250813 334516 250873
rect 334550 250813 334556 250873
rect 334505 250801 334556 250813
rect 334668 250873 334727 250885
rect 334668 250813 334674 250873
rect 334708 250813 334727 250873
rect 334668 250801 334727 250813
rect 334771 250885 334805 251061
rect 334842 250957 334934 250963
rect 334842 250923 334854 250957
rect 334922 250923 334934 250957
rect 334842 250917 334934 250923
rect 335118 250957 335210 250963
rect 335118 250923 335130 250957
rect 335198 250923 335210 250957
rect 335118 250917 335210 250923
rect 334969 250885 334999 250909
rect 334771 250873 334832 250885
rect 334771 250813 334792 250873
rect 334826 250813 334832 250873
rect 334771 250801 334832 250813
rect 334944 250873 334999 250885
rect 334944 250813 334950 250873
rect 334984 250813 334999 250873
rect 334944 250801 334999 250813
rect 334505 250637 334535 250801
rect 334693 250799 334727 250801
rect 334566 250763 334658 250769
rect 334566 250729 334578 250763
rect 334646 250729 334658 250763
rect 334566 250723 334658 250729
rect 334842 250763 334934 250769
rect 334842 250729 334854 250763
rect 334922 250729 334934 250763
rect 334842 250723 334934 250729
rect 334969 250637 334999 250801
rect 335055 250885 335085 250913
rect 335243 250885 335277 251061
rect 335055 250873 335108 250885
rect 335055 250813 335068 250873
rect 335102 250813 335108 250873
rect 335055 250801 335108 250813
rect 335220 250873 335277 250885
rect 335220 250813 335226 250873
rect 335260 250813 335277 250873
rect 335220 250801 335277 250813
rect 335055 250637 335085 250801
rect 335243 250797 335277 250801
rect 335327 250885 335361 251061
rect 335394 250957 335486 250963
rect 335394 250923 335406 250957
rect 335474 250923 335486 250957
rect 335394 250917 335486 250923
rect 335670 250957 335762 250963
rect 335670 250923 335682 250957
rect 335750 250923 335762 250957
rect 335670 250917 335762 250923
rect 335515 250885 335545 250899
rect 335327 250873 335384 250885
rect 335327 250813 335344 250873
rect 335378 250813 335384 250873
rect 335327 250801 335384 250813
rect 335496 250873 335545 250885
rect 335496 250813 335502 250873
rect 335536 250813 335545 250873
rect 335496 250801 335545 250813
rect 335327 250795 335361 250801
rect 335118 250763 335210 250769
rect 335118 250729 335130 250763
rect 335198 250729 335210 250763
rect 335118 250723 335210 250729
rect 335394 250763 335486 250769
rect 335394 250729 335406 250763
rect 335474 250729 335486 250763
rect 335394 250723 335486 250729
rect 335515 250637 335545 250801
rect 335607 250885 335637 250897
rect 335795 250885 335829 251061
rect 335607 250873 335660 250885
rect 335607 250813 335620 250873
rect 335654 250813 335660 250873
rect 335607 250801 335660 250813
rect 335772 250873 335829 250885
rect 335772 250813 335778 250873
rect 335812 250813 335829 250873
rect 335772 250801 335829 250813
rect 335607 250637 335637 250801
rect 335795 250797 335829 250801
rect 335879 250885 335913 251061
rect 335946 250957 336038 250963
rect 335946 250923 335958 250957
rect 336026 250923 336038 250957
rect 335946 250917 336038 250923
rect 336222 250957 336314 250963
rect 336222 250923 336234 250957
rect 336302 250923 336314 250957
rect 336222 250917 336314 250923
rect 336071 250885 336101 250899
rect 335879 250873 335936 250885
rect 335879 250813 335896 250873
rect 335930 250813 335936 250873
rect 335879 250801 335936 250813
rect 336048 250873 336101 250885
rect 336048 250813 336054 250873
rect 336088 250813 336101 250873
rect 336048 250801 336101 250813
rect 335879 250799 335913 250801
rect 335670 250763 335762 250769
rect 335670 250729 335682 250763
rect 335750 250729 335762 250763
rect 335670 250723 335762 250729
rect 335946 250763 336038 250769
rect 335946 250729 335958 250763
rect 336026 250729 336038 250763
rect 335946 250723 336038 250729
rect 336071 250637 336101 250801
rect 336155 250885 336185 250899
rect 336349 250885 336383 251061
rect 336155 250873 336212 250885
rect 336155 250813 336172 250873
rect 336206 250813 336212 250873
rect 336155 250801 336212 250813
rect 336324 250873 336383 250885
rect 336324 250813 336330 250873
rect 336364 250813 336383 250873
rect 336324 250803 336383 250813
rect 336427 250885 336461 251061
rect 336498 250957 336590 250963
rect 336498 250923 336510 250957
rect 336578 250923 336590 250957
rect 336498 250917 336590 250923
rect 336621 250885 336651 250899
rect 336427 250873 336488 250885
rect 336427 250813 336448 250873
rect 336482 250813 336488 250873
rect 336324 250801 336370 250803
rect 336427 250801 336488 250813
rect 336600 250873 336651 250885
rect 336600 250813 336606 250873
rect 336640 250813 336651 250873
rect 336600 250801 336651 250813
rect 336741 250809 336775 251061
rect 336155 250637 336185 250801
rect 336222 250763 336314 250769
rect 336222 250729 336234 250763
rect 336302 250729 336314 250763
rect 336222 250723 336314 250729
rect 336498 250763 336590 250769
rect 336498 250729 336510 250763
rect 336578 250729 336590 250763
rect 336498 250723 336590 250729
rect 336621 250637 336651 250801
rect 322484 250595 336653 250637
rect 336611 250593 336653 250595
rect 146202 250132 148512 250136
rect 148776 250132 150882 250136
rect 146202 249536 150882 250132
rect 60798 248220 60958 248820
rect 61558 248220 61758 248820
rect 60798 248060 61758 248220
rect 52310 239406 52640 240230
rect 53366 239406 53762 240230
rect 52310 238812 53762 239406
rect 141434 240026 142886 248942
rect 146202 248616 147162 249536
rect 146202 248016 146362 248616
rect 146962 248016 147162 248616
rect 146202 247856 147162 248016
rect 149922 248616 150882 249536
rect 233248 249098 233572 250500
rect 326663 250489 326803 250501
rect 326663 250433 326703 250489
rect 326781 250433 326803 250489
rect 326663 249819 326803 250433
rect 337591 250134 339092 251061
rect 323035 249619 326849 249819
rect 233250 248754 233514 249098
rect 149922 248016 150082 248616
rect 150682 248016 150882 248616
rect 149922 247856 150882 248016
rect 141434 239202 141764 240026
rect 142490 239202 142886 240026
rect 141434 238608 142886 239202
rect 232688 239838 234140 248754
rect 323035 247388 323235 249619
rect 411258 249730 412348 251411
rect 413127 251233 413169 251411
rect 413285 251409 413291 251411
rect 413325 251409 413331 251469
rect 413285 251397 413331 251409
rect 413443 251469 413506 251481
rect 413443 251409 413449 251469
rect 413483 251409 413506 251469
rect 413443 251397 413506 251409
rect 413466 251391 413506 251397
rect 413548 251481 413588 251657
rect 413617 251553 413709 251559
rect 413617 251519 413629 251553
rect 413697 251519 413709 251553
rect 413617 251513 413709 251519
rect 413893 251553 413985 251559
rect 413893 251519 413905 251553
rect 413973 251519 413985 251553
rect 413893 251513 413985 251519
rect 413742 251481 413772 251489
rect 413548 251469 413607 251481
rect 413548 251409 413567 251469
rect 413601 251409 413607 251469
rect 413548 251397 413607 251409
rect 413719 251469 413772 251481
rect 413719 251409 413725 251469
rect 413759 251409 413772 251469
rect 413719 251397 413772 251409
rect 413548 251393 413588 251397
rect 413341 251359 413433 251365
rect 413341 251325 413353 251359
rect 413421 251325 413433 251359
rect 413341 251319 413433 251325
rect 413617 251359 413709 251365
rect 413617 251325 413629 251359
rect 413697 251325 413709 251359
rect 413617 251319 413709 251325
rect 413742 251233 413772 251397
rect 413828 251481 413858 251489
rect 414024 251481 414064 251657
rect 413828 251469 413883 251481
rect 413828 251409 413843 251469
rect 413877 251409 413883 251469
rect 413828 251397 413883 251409
rect 413995 251469 414064 251481
rect 413995 251409 414001 251469
rect 414035 251409 414064 251469
rect 413995 251397 414064 251409
rect 413828 251233 413858 251397
rect 414024 251393 414064 251397
rect 414092 251481 414132 251657
rect 414169 251553 414261 251559
rect 414169 251519 414181 251553
rect 414249 251519 414261 251553
rect 414169 251513 414261 251519
rect 414445 251553 414537 251559
rect 414445 251519 414457 251553
rect 414525 251519 414537 251553
rect 414445 251513 414537 251519
rect 414296 251481 414326 251489
rect 414092 251469 414159 251481
rect 414092 251409 414119 251469
rect 414153 251409 414159 251469
rect 414092 251397 414159 251409
rect 414271 251469 414326 251481
rect 414271 251409 414277 251469
rect 414311 251409 414326 251469
rect 414271 251397 414326 251409
rect 414092 251393 414132 251397
rect 413893 251359 413985 251365
rect 413893 251325 413905 251359
rect 413973 251325 413985 251359
rect 413893 251319 413985 251325
rect 414169 251359 414261 251365
rect 414169 251325 414181 251359
rect 414249 251325 414261 251359
rect 414169 251319 414261 251325
rect 414296 251233 414326 251397
rect 414382 251481 414412 251489
rect 414572 251481 414612 251657
rect 414382 251469 414435 251481
rect 414382 251409 414395 251469
rect 414429 251409 414435 251469
rect 414382 251397 414435 251409
rect 414547 251469 414612 251481
rect 414547 251409 414553 251469
rect 414587 251409 414612 251469
rect 414547 251397 414612 251409
rect 414382 251233 414412 251397
rect 414572 251389 414612 251397
rect 414644 251481 414684 251657
rect 414721 251553 414813 251559
rect 414721 251519 414733 251553
rect 414801 251519 414813 251553
rect 414721 251513 414813 251519
rect 414997 251553 415089 251559
rect 414997 251519 415009 251553
rect 415077 251519 415089 251553
rect 414997 251513 415089 251519
rect 414844 251481 414874 251489
rect 414644 251469 414711 251481
rect 414644 251409 414671 251469
rect 414705 251409 414711 251469
rect 414644 251397 414711 251409
rect 414823 251469 414874 251481
rect 414823 251409 414829 251469
rect 414863 251409 414874 251469
rect 414823 251397 414874 251409
rect 414644 251393 414684 251397
rect 414445 251359 414537 251365
rect 414445 251325 414457 251359
rect 414525 251325 414537 251359
rect 414445 251319 414537 251325
rect 414721 251359 414813 251365
rect 414721 251325 414733 251359
rect 414801 251325 414813 251359
rect 414721 251319 414813 251325
rect 414844 251233 414874 251397
rect 414936 251481 414966 251487
rect 415124 251481 415164 251657
rect 414936 251469 414987 251481
rect 414936 251409 414947 251469
rect 414981 251409 414987 251469
rect 414936 251397 414987 251409
rect 415099 251469 415164 251481
rect 415099 251409 415105 251469
rect 415139 251409 415164 251469
rect 415099 251397 415164 251409
rect 415204 251481 415244 251657
rect 415273 251553 415365 251559
rect 415273 251519 415285 251553
rect 415353 251519 415365 251553
rect 415273 251513 415365 251519
rect 415549 251553 415641 251559
rect 415549 251519 415561 251553
rect 415629 251519 415641 251553
rect 415549 251513 415641 251519
rect 415394 251481 415424 251487
rect 415204 251469 415263 251481
rect 415204 251409 415223 251469
rect 415257 251409 415263 251469
rect 415204 251397 415263 251409
rect 415375 251469 415424 251481
rect 415375 251409 415381 251469
rect 415415 251409 415424 251469
rect 415375 251397 415424 251409
rect 414936 251233 414966 251397
rect 414997 251359 415089 251365
rect 414997 251325 415009 251359
rect 415077 251325 415089 251359
rect 414997 251319 415089 251325
rect 415273 251359 415365 251365
rect 415273 251325 415285 251359
rect 415353 251325 415365 251359
rect 415273 251319 415365 251325
rect 415394 251233 415424 251397
rect 415486 251481 415516 251485
rect 415678 251481 415718 251657
rect 415486 251469 415539 251481
rect 415486 251409 415499 251469
rect 415533 251409 415539 251469
rect 415486 251397 415539 251409
rect 415651 251469 415718 251481
rect 415651 251409 415657 251469
rect 415691 251409 415718 251469
rect 415651 251397 415718 251409
rect 415486 251233 415516 251397
rect 415678 251393 415718 251397
rect 415752 251481 415792 251657
rect 415825 251553 415917 251559
rect 415825 251519 415837 251553
rect 415905 251519 415917 251553
rect 415825 251513 415917 251519
rect 416101 251553 416193 251559
rect 416101 251519 416113 251553
rect 416181 251519 416193 251553
rect 416101 251513 416193 251519
rect 415950 251481 415980 251485
rect 415752 251469 415815 251481
rect 415752 251409 415775 251469
rect 415809 251409 415815 251469
rect 415752 251397 415815 251409
rect 415927 251469 415980 251481
rect 415927 251409 415933 251469
rect 415967 251409 415980 251469
rect 415927 251397 415980 251409
rect 415752 251395 415792 251397
rect 415549 251359 415641 251365
rect 415549 251325 415561 251359
rect 415629 251325 415641 251359
rect 415549 251319 415641 251325
rect 415825 251359 415917 251365
rect 415825 251325 415837 251359
rect 415905 251325 415917 251359
rect 415825 251319 415917 251325
rect 415950 251233 415980 251397
rect 416038 251481 416068 251483
rect 416230 251481 416270 251657
rect 416038 251469 416091 251481
rect 416038 251409 416051 251469
rect 416085 251409 416091 251469
rect 416038 251397 416091 251409
rect 416203 251469 416270 251481
rect 416203 251409 416209 251469
rect 416243 251409 416270 251469
rect 416203 251397 416270 251409
rect 416038 251233 416068 251397
rect 416230 251391 416270 251397
rect 416300 251481 416340 251657
rect 416377 251553 416469 251559
rect 416377 251519 416389 251553
rect 416457 251519 416469 251553
rect 416377 251513 416469 251519
rect 416653 251553 416745 251559
rect 416653 251519 416665 251553
rect 416733 251519 416745 251553
rect 416653 251513 416745 251519
rect 416500 251481 416530 251483
rect 416300 251469 416367 251481
rect 416300 251409 416327 251469
rect 416361 251409 416367 251469
rect 416300 251397 416367 251409
rect 416479 251469 416530 251481
rect 416479 251409 416485 251469
rect 416519 251409 416530 251469
rect 416479 251397 416530 251409
rect 416300 251395 416340 251397
rect 416101 251359 416193 251365
rect 416377 251363 416469 251365
rect 416101 251325 416113 251359
rect 416181 251325 416193 251359
rect 416374 251359 416469 251363
rect 416374 251330 416389 251359
rect 416101 251319 416193 251325
rect 416377 251325 416389 251330
rect 416457 251325 416469 251359
rect 416377 251319 416469 251325
rect 416500 251233 416530 251397
rect 416588 251481 416618 251483
rect 416778 251481 416818 251657
rect 416588 251469 416643 251481
rect 416588 251409 416603 251469
rect 416637 251409 416643 251469
rect 416588 251397 416643 251409
rect 416755 251469 416818 251481
rect 416755 251409 416761 251469
rect 416795 251409 416818 251469
rect 416755 251397 416818 251409
rect 416588 251233 416618 251397
rect 416778 251391 416818 251397
rect 416856 251481 416896 251657
rect 416929 251553 417021 251559
rect 416929 251519 416941 251553
rect 417009 251519 417021 251553
rect 416929 251513 417021 251519
rect 417205 251553 417297 251559
rect 417205 251519 417217 251553
rect 417285 251519 417297 251553
rect 417205 251513 417297 251519
rect 417052 251481 417082 251485
rect 416856 251469 416919 251481
rect 416856 251409 416879 251469
rect 416913 251409 416919 251469
rect 416856 251397 416919 251409
rect 417031 251469 417082 251481
rect 417031 251409 417037 251469
rect 417071 251409 417082 251469
rect 417031 251397 417082 251409
rect 416856 251395 416896 251397
rect 416653 251359 416745 251365
rect 416653 251325 416665 251359
rect 416733 251325 416745 251359
rect 416653 251319 416745 251325
rect 416929 251359 417021 251365
rect 416929 251325 416941 251359
rect 417009 251325 417021 251359
rect 416929 251319 417021 251325
rect 417052 251233 417082 251397
rect 417140 251481 417170 251485
rect 417332 251481 417372 251657
rect 417140 251469 417195 251481
rect 417140 251409 417155 251469
rect 417189 251409 417195 251469
rect 417140 251397 417195 251409
rect 417307 251469 417372 251481
rect 417307 251409 417313 251469
rect 417347 251409 417372 251469
rect 417307 251397 417372 251409
rect 417140 251233 417170 251397
rect 417332 251383 417372 251397
rect 417410 251481 417450 251657
rect 417481 251553 417573 251559
rect 417481 251519 417493 251553
rect 417561 251519 417573 251553
rect 417481 251513 417573 251519
rect 417757 251553 417849 251559
rect 417757 251519 417769 251553
rect 417837 251519 417849 251553
rect 417757 251513 417849 251519
rect 417604 251481 417634 251485
rect 417410 251469 417471 251481
rect 417410 251409 417431 251469
rect 417465 251409 417471 251469
rect 417410 251397 417471 251409
rect 417583 251469 417634 251481
rect 417583 251409 417589 251469
rect 417623 251409 417634 251469
rect 417583 251397 417634 251409
rect 417410 251391 417450 251397
rect 417205 251359 417297 251365
rect 417205 251325 417217 251359
rect 417285 251325 417297 251359
rect 417205 251319 417297 251325
rect 417481 251359 417573 251365
rect 417481 251325 417493 251359
rect 417561 251325 417573 251359
rect 417481 251319 417573 251325
rect 417604 251233 417634 251397
rect 417696 251481 417726 251485
rect 417888 251481 417928 251657
rect 417696 251469 417747 251481
rect 417696 251409 417707 251469
rect 417741 251409 417747 251469
rect 417696 251397 417747 251409
rect 417859 251469 417928 251481
rect 417859 251409 417865 251469
rect 417899 251409 417928 251469
rect 417859 251397 417928 251409
rect 417962 251481 418002 251657
rect 418033 251553 418125 251559
rect 418033 251519 418045 251553
rect 418113 251519 418125 251553
rect 418033 251513 418125 251519
rect 418309 251553 418401 251559
rect 418309 251519 418321 251553
rect 418389 251519 418401 251553
rect 418309 251513 418401 251519
rect 418158 251481 418188 251495
rect 417962 251469 418023 251481
rect 417962 251409 417983 251469
rect 418017 251409 418023 251469
rect 417962 251397 418023 251409
rect 418135 251469 418188 251481
rect 418135 251409 418141 251469
rect 418175 251409 418188 251469
rect 418135 251397 418188 251409
rect 417696 251233 417726 251397
rect 417888 251393 417928 251397
rect 417757 251359 417849 251365
rect 417757 251325 417769 251359
rect 417837 251325 417849 251359
rect 417757 251319 417849 251325
rect 418033 251359 418125 251365
rect 418033 251325 418045 251359
rect 418113 251325 418125 251359
rect 418033 251319 418125 251325
rect 418158 251233 418188 251397
rect 418244 251481 418274 251493
rect 418432 251481 418466 251657
rect 418244 251469 418299 251481
rect 418244 251409 418259 251469
rect 418293 251409 418299 251469
rect 418244 251397 418299 251409
rect 418411 251469 418466 251481
rect 418411 251409 418417 251469
rect 418451 251409 418466 251469
rect 418411 251397 418466 251409
rect 418244 251233 418274 251397
rect 418432 251393 418466 251397
rect 418522 251481 418556 251657
rect 418585 251553 418677 251559
rect 418585 251519 418597 251553
rect 418665 251519 418677 251553
rect 418585 251513 418677 251519
rect 418861 251553 418953 251559
rect 418861 251519 418873 251553
rect 418941 251519 418953 251553
rect 418861 251513 418953 251519
rect 418712 251481 418742 251491
rect 418522 251469 418575 251481
rect 418522 251409 418535 251469
rect 418569 251409 418575 251469
rect 418522 251397 418575 251409
rect 418687 251469 418742 251481
rect 418687 251409 418693 251469
rect 418727 251409 418742 251469
rect 418687 251397 418742 251409
rect 418522 251393 418556 251397
rect 418309 251359 418401 251365
rect 418309 251325 418321 251359
rect 418389 251325 418401 251359
rect 418309 251319 418401 251325
rect 418585 251359 418677 251365
rect 418585 251325 418597 251359
rect 418665 251325 418677 251359
rect 418585 251319 418677 251325
rect 418712 251233 418742 251397
rect 418798 251481 418828 251491
rect 418988 251481 419022 251657
rect 418798 251469 418851 251481
rect 418798 251409 418811 251469
rect 418845 251409 418851 251469
rect 418798 251397 418851 251409
rect 418963 251469 419022 251481
rect 418963 251409 418969 251469
rect 419003 251409 419022 251469
rect 418963 251397 419022 251409
rect 419072 251481 419106 251657
rect 419137 251553 419229 251559
rect 419137 251519 419149 251553
rect 419217 251519 419229 251553
rect 419137 251513 419229 251519
rect 419264 251481 419298 251495
rect 419072 251469 419127 251481
rect 419072 251409 419087 251469
rect 419121 251409 419127 251469
rect 419072 251397 419127 251409
rect 419239 251469 419298 251481
rect 419239 251409 419245 251469
rect 419279 251409 419298 251469
rect 419239 251397 419298 251409
rect 418798 251233 418828 251397
rect 418988 251393 419022 251397
rect 418861 251359 418953 251365
rect 418861 251325 418873 251359
rect 418941 251325 418953 251359
rect 418861 251319 418953 251325
rect 419137 251359 419229 251365
rect 419137 251325 419149 251359
rect 419217 251325 419229 251359
rect 419137 251319 419229 251325
rect 419264 251233 419298 251397
rect 419346 251481 419380 251657
rect 419413 251553 419505 251559
rect 419413 251519 419425 251553
rect 419493 251519 419505 251553
rect 419413 251513 419505 251519
rect 419689 251553 419781 251559
rect 419689 251519 419701 251553
rect 419769 251519 419781 251553
rect 419689 251513 419781 251519
rect 419538 251481 419568 251493
rect 419346 251469 419403 251481
rect 419346 251409 419363 251469
rect 419397 251409 419403 251469
rect 419346 251397 419403 251409
rect 419515 251469 419568 251481
rect 419515 251409 419521 251469
rect 419555 251409 419568 251469
rect 419515 251397 419568 251409
rect 419346 251395 419380 251397
rect 419413 251359 419505 251365
rect 419413 251325 419425 251359
rect 419493 251325 419505 251359
rect 419413 251319 419505 251325
rect 419538 251233 419568 251397
rect 419626 251481 419656 251495
rect 419816 251481 419850 251657
rect 419626 251469 419679 251481
rect 419626 251409 419639 251469
rect 419673 251409 419679 251469
rect 419626 251397 419679 251409
rect 419791 251469 419850 251481
rect 419791 251409 419797 251469
rect 419831 251409 419850 251469
rect 419791 251397 419850 251409
rect 419902 251481 419936 251657
rect 419974 251595 420189 251605
rect 419974 251559 420104 251595
rect 419965 251553 420104 251559
rect 419965 251519 419977 251553
rect 420045 251535 420104 251553
rect 420164 251535 420189 251595
rect 420045 251525 420189 251535
rect 420241 251553 420333 251559
rect 420045 251519 420057 251525
rect 419965 251513 420057 251519
rect 420241 251519 420253 251553
rect 420321 251519 420333 251553
rect 420241 251513 420333 251519
rect 420086 251481 420116 251495
rect 419902 251469 419955 251481
rect 419902 251409 419915 251469
rect 419949 251409 419955 251469
rect 419902 251397 419955 251409
rect 420067 251469 420116 251481
rect 420067 251409 420073 251469
rect 420107 251409 420116 251469
rect 420067 251397 420116 251409
rect 419626 251233 419656 251397
rect 419902 251391 419936 251397
rect 419689 251359 419781 251365
rect 419689 251325 419701 251359
rect 419769 251325 419781 251359
rect 419965 251359 420057 251365
rect 419965 251340 419977 251359
rect 419689 251319 419781 251325
rect 419829 251335 419977 251340
rect 419829 251280 419839 251335
rect 419904 251325 419977 251335
rect 420045 251325 420057 251359
rect 419904 251319 420057 251325
rect 419904 251290 420044 251319
rect 419904 251280 419914 251290
rect 419829 251275 419914 251280
rect 420086 251233 420116 251397
rect 420178 251481 420208 251495
rect 420368 251481 420402 251657
rect 420178 251469 420231 251481
rect 420178 251409 420191 251469
rect 420225 251409 420231 251469
rect 420178 251397 420231 251409
rect 420343 251469 420402 251481
rect 420343 251409 420349 251469
rect 420383 251409 420402 251469
rect 420343 251399 420402 251409
rect 420454 251481 420488 251657
rect 420517 251553 420609 251559
rect 420517 251519 420529 251553
rect 420597 251519 420609 251553
rect 420517 251513 420609 251519
rect 420793 251553 420885 251559
rect 420793 251519 420805 251553
rect 420873 251519 420885 251553
rect 420793 251513 420885 251519
rect 420640 251481 420670 251495
rect 420454 251469 420507 251481
rect 420454 251409 420467 251469
rect 420501 251409 420507 251469
rect 420343 251397 420389 251399
rect 420454 251397 420507 251409
rect 420619 251469 420670 251481
rect 420619 251409 420625 251469
rect 420659 251409 420670 251469
rect 420619 251397 420670 251409
rect 420178 251233 420208 251397
rect 420454 251395 420488 251397
rect 420241 251359 420333 251365
rect 420241 251325 420253 251359
rect 420321 251325 420333 251359
rect 420241 251319 420333 251325
rect 420517 251359 420609 251365
rect 420517 251325 420529 251359
rect 420597 251325 420609 251359
rect 420517 251319 420609 251325
rect 420640 251233 420670 251397
rect 420732 251481 420762 251495
rect 420918 251481 420952 251657
rect 420732 251469 420783 251481
rect 420732 251409 420743 251469
rect 420777 251409 420783 251469
rect 420732 251397 420783 251409
rect 420895 251469 420952 251481
rect 420895 251409 420901 251469
rect 420935 251409 420952 251469
rect 420895 251397 420952 251409
rect 420732 251233 420762 251397
rect 420918 251395 420952 251397
rect 421006 251481 421040 251657
rect 421069 251553 421161 251559
rect 421069 251519 421081 251553
rect 421149 251519 421161 251553
rect 421069 251513 421161 251519
rect 421345 251553 421437 251559
rect 421345 251519 421357 251553
rect 421425 251519 421437 251553
rect 421345 251513 421437 251519
rect 421192 251481 421222 251495
rect 421006 251469 421059 251481
rect 421006 251409 421019 251469
rect 421053 251409 421059 251469
rect 421006 251397 421059 251409
rect 421171 251469 421222 251481
rect 421171 251409 421177 251469
rect 421211 251409 421222 251469
rect 421171 251397 421222 251409
rect 421006 251393 421040 251397
rect 420793 251359 420885 251365
rect 420793 251325 420805 251359
rect 420873 251325 420885 251359
rect 420793 251319 420885 251325
rect 421069 251359 421161 251365
rect 421069 251325 421081 251359
rect 421149 251325 421161 251359
rect 421069 251319 421161 251325
rect 421192 251233 421222 251397
rect 421278 251481 421308 251495
rect 421474 251481 421508 251657
rect 421278 251469 421335 251481
rect 421278 251409 421295 251469
rect 421329 251409 421335 251469
rect 421278 251397 421335 251409
rect 421447 251469 421508 251481
rect 421447 251409 421453 251469
rect 421487 251409 421508 251469
rect 421447 251397 421508 251409
rect 421278 251233 421308 251397
rect 421474 251389 421508 251397
rect 421556 251481 421590 251657
rect 421621 251553 421713 251559
rect 421621 251519 421633 251553
rect 421701 251519 421713 251553
rect 421621 251513 421713 251519
rect 421897 251553 421989 251559
rect 421897 251519 421909 251553
rect 421977 251519 421989 251553
rect 421897 251513 421989 251519
rect 421746 251481 421776 251495
rect 421556 251469 421611 251481
rect 421556 251409 421571 251469
rect 421605 251409 421611 251469
rect 421556 251397 421611 251409
rect 421723 251469 421776 251481
rect 421723 251409 421729 251469
rect 421763 251409 421776 251469
rect 421723 251397 421776 251409
rect 421556 251395 421590 251397
rect 421345 251359 421437 251365
rect 421345 251325 421357 251359
rect 421425 251325 421437 251359
rect 421345 251319 421437 251325
rect 421621 251359 421713 251365
rect 421621 251325 421633 251359
rect 421701 251325 421713 251359
rect 421621 251319 421713 251325
rect 421746 251233 421776 251397
rect 421834 251481 421864 251493
rect 422028 251481 422062 251657
rect 421834 251469 421887 251481
rect 421834 251409 421847 251469
rect 421881 251409 421887 251469
rect 421834 251397 421887 251409
rect 421999 251469 422062 251481
rect 421999 251409 422005 251469
rect 422039 251409 422062 251469
rect 421999 251397 422062 251409
rect 421834 251233 421864 251397
rect 422028 251393 422062 251397
rect 422106 251481 422140 251657
rect 422173 251553 422265 251559
rect 422173 251519 422185 251553
rect 422253 251519 422265 251553
rect 422173 251513 422265 251519
rect 422449 251553 422541 251559
rect 422449 251519 422461 251553
rect 422529 251519 422541 251553
rect 422449 251513 422541 251519
rect 422298 251481 422328 251497
rect 422106 251469 422163 251481
rect 422106 251409 422123 251469
rect 422157 251409 422163 251469
rect 422106 251397 422163 251409
rect 422275 251469 422328 251481
rect 422275 251409 422281 251469
rect 422315 251409 422328 251469
rect 422275 251397 422328 251409
rect 422106 251395 422140 251397
rect 421897 251359 421989 251365
rect 421897 251325 421909 251359
rect 421977 251325 421989 251359
rect 421897 251319 421989 251325
rect 422173 251359 422265 251365
rect 422173 251325 422185 251359
rect 422253 251325 422265 251359
rect 422173 251319 422265 251325
rect 422298 251233 422328 251397
rect 422386 251481 422416 251497
rect 422584 251481 422618 251657
rect 422386 251469 422439 251481
rect 422386 251409 422399 251469
rect 422433 251409 422439 251469
rect 422386 251397 422439 251409
rect 422551 251469 422618 251481
rect 422551 251409 422557 251469
rect 422591 251409 422618 251469
rect 422551 251397 422618 251409
rect 422386 251233 422416 251397
rect 422584 251385 422618 251397
rect 422658 251481 422692 251657
rect 422725 251553 422817 251559
rect 422725 251519 422737 251553
rect 422805 251519 422817 251553
rect 422725 251513 422817 251519
rect 423001 251553 423093 251559
rect 423001 251519 423013 251553
rect 423081 251519 423093 251553
rect 423001 251513 423093 251519
rect 422848 251481 422878 251499
rect 422658 251469 422715 251481
rect 422658 251409 422675 251469
rect 422709 251409 422715 251469
rect 422658 251397 422715 251409
rect 422827 251469 422878 251481
rect 422827 251409 422833 251469
rect 422867 251409 422878 251469
rect 422827 251397 422878 251409
rect 422658 251389 422692 251397
rect 422449 251359 422541 251365
rect 422449 251325 422461 251359
rect 422529 251325 422541 251359
rect 422449 251319 422541 251325
rect 422725 251359 422817 251365
rect 422725 251325 422737 251359
rect 422805 251325 422817 251359
rect 422725 251319 422817 251325
rect 422848 251233 422878 251397
rect 422936 251481 422966 251497
rect 423128 251481 423162 251657
rect 422936 251469 422991 251481
rect 422936 251409 422951 251469
rect 422985 251409 422991 251469
rect 422936 251397 422991 251409
rect 423103 251469 423162 251481
rect 423103 251409 423109 251469
rect 423143 251409 423162 251469
rect 423103 251397 423162 251409
rect 422936 251233 422966 251397
rect 423128 251385 423162 251397
rect 423208 251481 423242 251657
rect 423277 251553 423369 251559
rect 423277 251519 423289 251553
rect 423357 251519 423369 251553
rect 423277 251513 423369 251519
rect 423553 251553 423645 251559
rect 423553 251519 423565 251553
rect 423633 251519 423645 251553
rect 423553 251513 423645 251519
rect 423400 251481 423430 251497
rect 423208 251469 423267 251481
rect 423208 251409 423227 251469
rect 423261 251409 423267 251469
rect 423208 251397 423267 251409
rect 423379 251469 423430 251481
rect 423379 251409 423385 251469
rect 423419 251409 423430 251469
rect 423379 251397 423430 251409
rect 423208 251383 423242 251397
rect 423001 251359 423093 251365
rect 423001 251325 423013 251359
rect 423081 251325 423093 251359
rect 423001 251319 423093 251325
rect 423277 251359 423369 251365
rect 423277 251325 423289 251359
rect 423357 251325 423369 251359
rect 423277 251319 423369 251325
rect 423400 251233 423430 251397
rect 423488 251481 423518 251499
rect 423684 251481 423718 251657
rect 423488 251469 423543 251481
rect 423488 251409 423503 251469
rect 423537 251409 423543 251469
rect 423488 251397 423543 251409
rect 423655 251469 423718 251481
rect 423655 251409 423661 251469
rect 423695 251409 423718 251469
rect 423655 251397 423718 251409
rect 423488 251233 423518 251397
rect 423684 251385 423718 251397
rect 423758 251481 423792 251657
rect 423829 251553 423921 251559
rect 423829 251519 423841 251553
rect 423909 251519 423921 251553
rect 423829 251513 423921 251519
rect 424105 251553 424197 251559
rect 424105 251519 424117 251553
rect 424185 251519 424197 251553
rect 424105 251513 424197 251519
rect 423952 251481 423982 251497
rect 423758 251469 423819 251481
rect 423758 251409 423779 251469
rect 423813 251409 423819 251469
rect 423758 251397 423819 251409
rect 423931 251469 423982 251481
rect 423931 251409 423937 251469
rect 423971 251409 423982 251469
rect 423931 251397 423982 251409
rect 423758 251383 423792 251397
rect 423553 251359 423645 251365
rect 423553 251325 423565 251359
rect 423633 251325 423645 251359
rect 423553 251319 423645 251325
rect 423829 251359 423921 251365
rect 423829 251325 423841 251359
rect 423909 251325 423921 251359
rect 423829 251319 423921 251325
rect 423952 251233 423982 251397
rect 424042 251481 424072 251499
rect 424234 251481 424268 251657
rect 424042 251469 424095 251481
rect 424042 251409 424055 251469
rect 424089 251409 424095 251469
rect 424042 251397 424095 251409
rect 424207 251469 424268 251481
rect 424207 251409 424213 251469
rect 424247 251409 424268 251469
rect 424207 251397 424268 251409
rect 424042 251233 424072 251397
rect 424234 251387 424268 251397
rect 424310 251481 424344 251657
rect 424381 251553 424473 251559
rect 424381 251519 424393 251553
rect 424461 251519 424473 251553
rect 424381 251513 424473 251519
rect 424657 251553 424749 251559
rect 424657 251519 424669 251553
rect 424737 251519 424749 251553
rect 424657 251513 424749 251519
rect 424504 251481 424534 251497
rect 424310 251469 424371 251481
rect 424310 251409 424331 251469
rect 424365 251409 424371 251469
rect 424310 251397 424371 251409
rect 424483 251469 424534 251481
rect 424483 251409 424489 251469
rect 424523 251409 424534 251469
rect 424483 251397 424534 251409
rect 424310 251387 424344 251397
rect 424105 251359 424197 251365
rect 424105 251325 424117 251359
rect 424185 251325 424197 251359
rect 424105 251319 424197 251325
rect 424381 251359 424473 251365
rect 424381 251325 424393 251359
rect 424461 251325 424473 251359
rect 424381 251319 424473 251325
rect 424504 251233 424534 251397
rect 424594 251481 424624 251499
rect 424784 251481 424818 251657
rect 424594 251469 424647 251481
rect 424594 251409 424607 251469
rect 424641 251409 424647 251469
rect 424594 251397 424647 251409
rect 424759 251469 424818 251481
rect 424759 251409 424765 251469
rect 424799 251409 424818 251469
rect 424759 251397 424818 251409
rect 424594 251233 424624 251397
rect 424784 251391 424818 251397
rect 424866 251481 424900 251657
rect 424933 251553 425025 251559
rect 424933 251519 424945 251553
rect 425013 251519 425025 251553
rect 424933 251513 425025 251519
rect 425209 251553 425301 251559
rect 425209 251519 425221 251553
rect 425289 251519 425301 251553
rect 425209 251513 425301 251519
rect 425058 251481 425088 251503
rect 424866 251469 424923 251481
rect 424866 251409 424883 251469
rect 424917 251409 424923 251469
rect 424866 251397 424923 251409
rect 425035 251469 425088 251481
rect 425035 251409 425041 251469
rect 425075 251409 425088 251469
rect 425035 251397 425088 251409
rect 424866 251389 424900 251397
rect 424657 251359 424749 251365
rect 424657 251325 424669 251359
rect 424737 251325 424749 251359
rect 424657 251319 424749 251325
rect 424933 251359 425025 251365
rect 424933 251325 424945 251359
rect 425013 251325 425025 251359
rect 424933 251319 425025 251325
rect 425058 251233 425088 251397
rect 425148 251481 425178 251505
rect 425336 251481 425370 251657
rect 425148 251469 425199 251481
rect 425148 251409 425159 251469
rect 425193 251409 425199 251469
rect 425148 251397 425199 251409
rect 425311 251469 425370 251481
rect 425311 251409 425317 251469
rect 425351 251409 425370 251469
rect 425311 251397 425370 251409
rect 425414 251481 425448 251657
rect 425485 251553 425577 251559
rect 425485 251519 425497 251553
rect 425565 251519 425577 251553
rect 425485 251513 425577 251519
rect 425761 251553 425853 251559
rect 425761 251519 425773 251553
rect 425841 251519 425853 251553
rect 425761 251513 425853 251519
rect 425612 251481 425642 251505
rect 425414 251469 425475 251481
rect 425414 251409 425435 251469
rect 425469 251409 425475 251469
rect 425414 251397 425475 251409
rect 425587 251469 425642 251481
rect 425587 251409 425593 251469
rect 425627 251409 425642 251469
rect 425587 251397 425642 251409
rect 425148 251233 425178 251397
rect 425336 251395 425370 251397
rect 425209 251359 425301 251365
rect 425209 251325 425221 251359
rect 425289 251325 425301 251359
rect 425209 251319 425301 251325
rect 425485 251359 425577 251365
rect 425485 251325 425497 251359
rect 425565 251325 425577 251359
rect 425485 251319 425577 251325
rect 425612 251233 425642 251397
rect 425698 251481 425728 251509
rect 425886 251481 425920 251657
rect 425698 251469 425751 251481
rect 425698 251409 425711 251469
rect 425745 251409 425751 251469
rect 425698 251397 425751 251409
rect 425863 251469 425920 251481
rect 425863 251409 425869 251469
rect 425903 251409 425920 251469
rect 425863 251397 425920 251409
rect 425698 251233 425728 251397
rect 425886 251393 425920 251397
rect 425970 251481 426004 251657
rect 426037 251553 426129 251559
rect 426037 251519 426049 251553
rect 426117 251519 426129 251553
rect 426037 251513 426129 251519
rect 426313 251553 426405 251559
rect 426313 251519 426325 251553
rect 426393 251519 426405 251553
rect 426313 251513 426405 251519
rect 426158 251481 426188 251495
rect 425970 251469 426027 251481
rect 425970 251409 425987 251469
rect 426021 251409 426027 251469
rect 425970 251397 426027 251409
rect 426139 251469 426188 251481
rect 426139 251409 426145 251469
rect 426179 251409 426188 251469
rect 426139 251397 426188 251409
rect 425970 251391 426004 251397
rect 425761 251359 425853 251365
rect 425761 251325 425773 251359
rect 425841 251325 425853 251359
rect 425761 251319 425853 251325
rect 426037 251359 426129 251365
rect 426037 251325 426049 251359
rect 426117 251325 426129 251359
rect 426037 251319 426129 251325
rect 426158 251233 426188 251397
rect 426250 251481 426280 251493
rect 426438 251481 426472 251657
rect 426250 251469 426303 251481
rect 426250 251409 426263 251469
rect 426297 251409 426303 251469
rect 426250 251397 426303 251409
rect 426415 251469 426472 251481
rect 426415 251409 426421 251469
rect 426455 251409 426472 251469
rect 426415 251397 426472 251409
rect 426250 251233 426280 251397
rect 426438 251393 426472 251397
rect 426522 251481 426556 251657
rect 426589 251553 426681 251559
rect 426589 251519 426601 251553
rect 426669 251519 426681 251553
rect 426589 251513 426681 251519
rect 426865 251553 426957 251559
rect 426865 251519 426877 251553
rect 426945 251519 426957 251553
rect 426865 251513 426957 251519
rect 426714 251481 426744 251495
rect 426522 251469 426579 251481
rect 426522 251409 426539 251469
rect 426573 251409 426579 251469
rect 426522 251397 426579 251409
rect 426691 251469 426744 251481
rect 426691 251409 426697 251469
rect 426731 251409 426744 251469
rect 426691 251397 426744 251409
rect 426522 251395 426556 251397
rect 426313 251359 426405 251365
rect 426313 251325 426325 251359
rect 426393 251325 426405 251359
rect 426313 251319 426405 251325
rect 426589 251359 426681 251365
rect 426589 251325 426601 251359
rect 426669 251325 426681 251359
rect 426589 251319 426681 251325
rect 426714 251233 426744 251397
rect 426798 251481 426828 251495
rect 426992 251481 427026 251657
rect 426798 251469 426855 251481
rect 426798 251409 426815 251469
rect 426849 251409 426855 251469
rect 426798 251397 426855 251409
rect 426967 251469 427026 251481
rect 426967 251409 426973 251469
rect 427007 251409 427026 251469
rect 426967 251399 427026 251409
rect 427070 251481 427104 251657
rect 427141 251553 427233 251559
rect 427141 251519 427153 251553
rect 427221 251519 427233 251553
rect 427141 251513 427233 251519
rect 427264 251481 427294 251495
rect 427070 251469 427131 251481
rect 427070 251409 427091 251469
rect 427125 251409 427131 251469
rect 426967 251397 427013 251399
rect 427070 251397 427131 251409
rect 427243 251469 427294 251481
rect 427243 251409 427249 251469
rect 427283 251409 427294 251469
rect 427243 251397 427294 251409
rect 427384 251405 427418 251657
rect 426798 251233 426828 251397
rect 426865 251359 426957 251365
rect 426865 251325 426877 251359
rect 426945 251325 426957 251359
rect 426865 251319 426957 251325
rect 427141 251359 427233 251365
rect 427141 251325 427153 251359
rect 427221 251325 427233 251359
rect 427141 251319 427233 251325
rect 427264 251233 427294 251397
rect 413127 251191 427296 251233
rect 427254 251189 427296 251191
rect 417306 251085 417446 251097
rect 417306 251029 417346 251085
rect 417424 251029 417446 251085
rect 417306 250415 417446 251029
rect 428318 250600 429188 251657
rect 411258 248634 412348 248640
rect 413138 250215 417492 250415
rect 337591 248627 339092 248633
rect 232688 239014 233018 239838
rect 233744 239014 234140 239838
rect 232688 238420 234140 239014
rect 322310 240230 323762 247388
rect 413138 245815 413338 250215
rect 428318 249724 429188 249730
rect 501258 251469 502348 252005
rect 518318 251723 519188 251755
rect 503461 251657 519188 251723
rect 503341 251553 503433 251559
rect 503341 251519 503353 251553
rect 503421 251519 503433 251553
rect 503341 251513 503433 251519
rect 503466 251481 503506 251657
rect 503285 251469 503331 251481
rect 501258 251411 503291 251469
rect 501258 249730 502348 251411
rect 503127 251233 503169 251411
rect 503285 251409 503291 251411
rect 503325 251409 503331 251469
rect 503285 251397 503331 251409
rect 503443 251469 503506 251481
rect 503443 251409 503449 251469
rect 503483 251409 503506 251469
rect 503443 251397 503506 251409
rect 503466 251391 503506 251397
rect 503548 251481 503588 251657
rect 503617 251553 503709 251559
rect 503617 251519 503629 251553
rect 503697 251519 503709 251553
rect 503617 251513 503709 251519
rect 503893 251553 503985 251559
rect 503893 251519 503905 251553
rect 503973 251519 503985 251553
rect 503893 251513 503985 251519
rect 503742 251481 503772 251489
rect 503548 251469 503607 251481
rect 503548 251409 503567 251469
rect 503601 251409 503607 251469
rect 503548 251397 503607 251409
rect 503719 251469 503772 251481
rect 503719 251409 503725 251469
rect 503759 251409 503772 251469
rect 503719 251397 503772 251409
rect 503548 251393 503588 251397
rect 503341 251359 503433 251365
rect 503341 251325 503353 251359
rect 503421 251325 503433 251359
rect 503341 251319 503433 251325
rect 503617 251359 503709 251365
rect 503617 251325 503629 251359
rect 503697 251325 503709 251359
rect 503617 251319 503709 251325
rect 503742 251233 503772 251397
rect 503828 251481 503858 251489
rect 504024 251481 504064 251657
rect 503828 251469 503883 251481
rect 503828 251409 503843 251469
rect 503877 251409 503883 251469
rect 503828 251397 503883 251409
rect 503995 251469 504064 251481
rect 503995 251409 504001 251469
rect 504035 251409 504064 251469
rect 503995 251397 504064 251409
rect 503828 251233 503858 251397
rect 504024 251393 504064 251397
rect 504092 251481 504132 251657
rect 504169 251553 504261 251559
rect 504169 251519 504181 251553
rect 504249 251519 504261 251553
rect 504169 251513 504261 251519
rect 504445 251553 504537 251559
rect 504445 251519 504457 251553
rect 504525 251519 504537 251553
rect 504445 251513 504537 251519
rect 504296 251481 504326 251489
rect 504092 251469 504159 251481
rect 504092 251409 504119 251469
rect 504153 251409 504159 251469
rect 504092 251397 504159 251409
rect 504271 251469 504326 251481
rect 504271 251409 504277 251469
rect 504311 251409 504326 251469
rect 504271 251397 504326 251409
rect 504092 251393 504132 251397
rect 503893 251359 503985 251365
rect 503893 251325 503905 251359
rect 503973 251325 503985 251359
rect 503893 251319 503985 251325
rect 504169 251359 504261 251365
rect 504169 251325 504181 251359
rect 504249 251325 504261 251359
rect 504169 251319 504261 251325
rect 504296 251233 504326 251397
rect 504382 251481 504412 251489
rect 504572 251481 504612 251657
rect 504382 251469 504435 251481
rect 504382 251409 504395 251469
rect 504429 251409 504435 251469
rect 504382 251397 504435 251409
rect 504547 251469 504612 251481
rect 504547 251409 504553 251469
rect 504587 251409 504612 251469
rect 504547 251397 504612 251409
rect 504382 251233 504412 251397
rect 504572 251389 504612 251397
rect 504644 251481 504684 251657
rect 504721 251553 504813 251559
rect 504721 251519 504733 251553
rect 504801 251519 504813 251553
rect 504721 251513 504813 251519
rect 504997 251553 505089 251559
rect 504997 251519 505009 251553
rect 505077 251519 505089 251553
rect 504997 251513 505089 251519
rect 504844 251481 504874 251489
rect 504644 251469 504711 251481
rect 504644 251409 504671 251469
rect 504705 251409 504711 251469
rect 504644 251397 504711 251409
rect 504823 251469 504874 251481
rect 504823 251409 504829 251469
rect 504863 251409 504874 251469
rect 504823 251397 504874 251409
rect 504644 251393 504684 251397
rect 504445 251359 504537 251365
rect 504445 251325 504457 251359
rect 504525 251325 504537 251359
rect 504445 251319 504537 251325
rect 504721 251359 504813 251365
rect 504721 251325 504733 251359
rect 504801 251325 504813 251359
rect 504721 251319 504813 251325
rect 504844 251233 504874 251397
rect 504936 251481 504966 251487
rect 505124 251481 505164 251657
rect 504936 251469 504987 251481
rect 504936 251409 504947 251469
rect 504981 251409 504987 251469
rect 504936 251397 504987 251409
rect 505099 251469 505164 251481
rect 505099 251409 505105 251469
rect 505139 251409 505164 251469
rect 505099 251397 505164 251409
rect 505204 251481 505244 251657
rect 505273 251553 505365 251559
rect 505273 251519 505285 251553
rect 505353 251519 505365 251553
rect 505273 251513 505365 251519
rect 505549 251553 505641 251559
rect 505549 251519 505561 251553
rect 505629 251519 505641 251553
rect 505549 251513 505641 251519
rect 505394 251481 505424 251487
rect 505204 251469 505263 251481
rect 505204 251409 505223 251469
rect 505257 251409 505263 251469
rect 505204 251397 505263 251409
rect 505375 251469 505424 251481
rect 505375 251409 505381 251469
rect 505415 251409 505424 251469
rect 505375 251397 505424 251409
rect 504936 251233 504966 251397
rect 504997 251359 505089 251365
rect 504997 251325 505009 251359
rect 505077 251325 505089 251359
rect 504997 251319 505089 251325
rect 505273 251359 505365 251365
rect 505273 251325 505285 251359
rect 505353 251325 505365 251359
rect 505273 251319 505365 251325
rect 505394 251233 505424 251397
rect 505486 251481 505516 251485
rect 505678 251481 505718 251657
rect 505486 251469 505539 251481
rect 505486 251409 505499 251469
rect 505533 251409 505539 251469
rect 505486 251397 505539 251409
rect 505651 251469 505718 251481
rect 505651 251409 505657 251469
rect 505691 251409 505718 251469
rect 505651 251397 505718 251409
rect 505486 251233 505516 251397
rect 505678 251393 505718 251397
rect 505752 251481 505792 251657
rect 505825 251553 505917 251559
rect 505825 251519 505837 251553
rect 505905 251519 505917 251553
rect 505825 251513 505917 251519
rect 506101 251553 506193 251559
rect 506101 251519 506113 251553
rect 506181 251519 506193 251553
rect 506101 251513 506193 251519
rect 505950 251481 505980 251485
rect 505752 251469 505815 251481
rect 505752 251409 505775 251469
rect 505809 251409 505815 251469
rect 505752 251397 505815 251409
rect 505927 251469 505980 251481
rect 505927 251409 505933 251469
rect 505967 251409 505980 251469
rect 505927 251397 505980 251409
rect 505752 251395 505792 251397
rect 505549 251359 505641 251365
rect 505549 251325 505561 251359
rect 505629 251325 505641 251359
rect 505549 251319 505641 251325
rect 505825 251359 505917 251365
rect 505825 251325 505837 251359
rect 505905 251325 505917 251359
rect 505825 251319 505917 251325
rect 505950 251233 505980 251397
rect 506038 251481 506068 251483
rect 506230 251481 506270 251657
rect 506038 251469 506091 251481
rect 506038 251409 506051 251469
rect 506085 251409 506091 251469
rect 506038 251397 506091 251409
rect 506203 251469 506270 251481
rect 506203 251409 506209 251469
rect 506243 251409 506270 251469
rect 506203 251397 506270 251409
rect 506038 251233 506068 251397
rect 506230 251391 506270 251397
rect 506300 251481 506340 251657
rect 506377 251553 506469 251559
rect 506377 251519 506389 251553
rect 506457 251519 506469 251553
rect 506377 251513 506469 251519
rect 506653 251553 506745 251559
rect 506653 251519 506665 251553
rect 506733 251519 506745 251553
rect 506653 251513 506745 251519
rect 506500 251481 506530 251483
rect 506300 251469 506367 251481
rect 506300 251409 506327 251469
rect 506361 251409 506367 251469
rect 506300 251397 506367 251409
rect 506479 251469 506530 251481
rect 506479 251409 506485 251469
rect 506519 251409 506530 251469
rect 506479 251397 506530 251409
rect 506300 251395 506340 251397
rect 506101 251359 506193 251365
rect 506377 251363 506469 251365
rect 506101 251325 506113 251359
rect 506181 251325 506193 251359
rect 506374 251359 506469 251363
rect 506374 251330 506389 251359
rect 506101 251319 506193 251325
rect 506377 251325 506389 251330
rect 506457 251325 506469 251359
rect 506377 251319 506469 251325
rect 506500 251233 506530 251397
rect 506588 251481 506618 251483
rect 506778 251481 506818 251657
rect 506588 251469 506643 251481
rect 506588 251409 506603 251469
rect 506637 251409 506643 251469
rect 506588 251397 506643 251409
rect 506755 251469 506818 251481
rect 506755 251409 506761 251469
rect 506795 251409 506818 251469
rect 506755 251397 506818 251409
rect 506588 251233 506618 251397
rect 506778 251391 506818 251397
rect 506856 251481 506896 251657
rect 506929 251553 507021 251559
rect 506929 251519 506941 251553
rect 507009 251519 507021 251553
rect 506929 251513 507021 251519
rect 507205 251553 507297 251559
rect 507205 251519 507217 251553
rect 507285 251519 507297 251553
rect 507205 251513 507297 251519
rect 507052 251481 507082 251485
rect 506856 251469 506919 251481
rect 506856 251409 506879 251469
rect 506913 251409 506919 251469
rect 506856 251397 506919 251409
rect 507031 251469 507082 251481
rect 507031 251409 507037 251469
rect 507071 251409 507082 251469
rect 507031 251397 507082 251409
rect 506856 251395 506896 251397
rect 506653 251359 506745 251365
rect 506653 251325 506665 251359
rect 506733 251325 506745 251359
rect 506653 251319 506745 251325
rect 506929 251359 507021 251365
rect 506929 251325 506941 251359
rect 507009 251325 507021 251359
rect 506929 251319 507021 251325
rect 507052 251233 507082 251397
rect 507140 251481 507170 251485
rect 507332 251481 507372 251657
rect 507140 251469 507195 251481
rect 507140 251409 507155 251469
rect 507189 251409 507195 251469
rect 507140 251397 507195 251409
rect 507307 251469 507372 251481
rect 507307 251409 507313 251469
rect 507347 251409 507372 251469
rect 507307 251397 507372 251409
rect 507140 251233 507170 251397
rect 507332 251383 507372 251397
rect 507410 251481 507450 251657
rect 507481 251553 507573 251559
rect 507481 251519 507493 251553
rect 507561 251519 507573 251553
rect 507481 251513 507573 251519
rect 507757 251553 507849 251559
rect 507757 251519 507769 251553
rect 507837 251519 507849 251553
rect 507757 251513 507849 251519
rect 507604 251481 507634 251485
rect 507410 251469 507471 251481
rect 507410 251409 507431 251469
rect 507465 251409 507471 251469
rect 507410 251397 507471 251409
rect 507583 251469 507634 251481
rect 507583 251409 507589 251469
rect 507623 251409 507634 251469
rect 507583 251397 507634 251409
rect 507410 251391 507450 251397
rect 507205 251359 507297 251365
rect 507205 251325 507217 251359
rect 507285 251325 507297 251359
rect 507205 251319 507297 251325
rect 507481 251359 507573 251365
rect 507481 251325 507493 251359
rect 507561 251325 507573 251359
rect 507481 251319 507573 251325
rect 507604 251233 507634 251397
rect 507696 251481 507726 251485
rect 507888 251481 507928 251657
rect 507696 251469 507747 251481
rect 507696 251409 507707 251469
rect 507741 251409 507747 251469
rect 507696 251397 507747 251409
rect 507859 251469 507928 251481
rect 507859 251409 507865 251469
rect 507899 251409 507928 251469
rect 507859 251397 507928 251409
rect 507962 251481 508002 251657
rect 508033 251553 508125 251559
rect 508033 251519 508045 251553
rect 508113 251519 508125 251553
rect 508033 251513 508125 251519
rect 508309 251553 508401 251559
rect 508309 251519 508321 251553
rect 508389 251519 508401 251553
rect 508309 251513 508401 251519
rect 508158 251481 508188 251495
rect 507962 251469 508023 251481
rect 507962 251409 507983 251469
rect 508017 251409 508023 251469
rect 507962 251397 508023 251409
rect 508135 251469 508188 251481
rect 508135 251409 508141 251469
rect 508175 251409 508188 251469
rect 508135 251397 508188 251409
rect 507696 251233 507726 251397
rect 507888 251393 507928 251397
rect 507757 251359 507849 251365
rect 507757 251325 507769 251359
rect 507837 251325 507849 251359
rect 507757 251319 507849 251325
rect 508033 251359 508125 251365
rect 508033 251325 508045 251359
rect 508113 251325 508125 251359
rect 508033 251319 508125 251325
rect 508158 251233 508188 251397
rect 508244 251481 508274 251493
rect 508432 251481 508466 251657
rect 508244 251469 508299 251481
rect 508244 251409 508259 251469
rect 508293 251409 508299 251469
rect 508244 251397 508299 251409
rect 508411 251469 508466 251481
rect 508411 251409 508417 251469
rect 508451 251409 508466 251469
rect 508411 251397 508466 251409
rect 508244 251233 508274 251397
rect 508432 251393 508466 251397
rect 508522 251481 508556 251657
rect 508585 251553 508677 251559
rect 508585 251519 508597 251553
rect 508665 251519 508677 251553
rect 508585 251513 508677 251519
rect 508861 251553 508953 251559
rect 508861 251519 508873 251553
rect 508941 251519 508953 251553
rect 508861 251513 508953 251519
rect 508712 251481 508742 251491
rect 508522 251469 508575 251481
rect 508522 251409 508535 251469
rect 508569 251409 508575 251469
rect 508522 251397 508575 251409
rect 508687 251469 508742 251481
rect 508687 251409 508693 251469
rect 508727 251409 508742 251469
rect 508687 251397 508742 251409
rect 508522 251393 508556 251397
rect 508309 251359 508401 251365
rect 508309 251325 508321 251359
rect 508389 251325 508401 251359
rect 508309 251319 508401 251325
rect 508585 251359 508677 251365
rect 508585 251325 508597 251359
rect 508665 251325 508677 251359
rect 508585 251319 508677 251325
rect 508712 251233 508742 251397
rect 508798 251481 508828 251491
rect 508988 251481 509022 251657
rect 508798 251469 508851 251481
rect 508798 251409 508811 251469
rect 508845 251409 508851 251469
rect 508798 251397 508851 251409
rect 508963 251469 509022 251481
rect 508963 251409 508969 251469
rect 509003 251409 509022 251469
rect 508963 251397 509022 251409
rect 509072 251481 509106 251657
rect 509137 251553 509229 251559
rect 509137 251519 509149 251553
rect 509217 251519 509229 251553
rect 509137 251513 509229 251519
rect 509264 251481 509298 251495
rect 509072 251469 509127 251481
rect 509072 251409 509087 251469
rect 509121 251409 509127 251469
rect 509072 251397 509127 251409
rect 509239 251469 509298 251481
rect 509239 251409 509245 251469
rect 509279 251409 509298 251469
rect 509239 251397 509298 251409
rect 508798 251233 508828 251397
rect 508988 251393 509022 251397
rect 508861 251359 508953 251365
rect 508861 251325 508873 251359
rect 508941 251325 508953 251359
rect 508861 251319 508953 251325
rect 509137 251359 509229 251365
rect 509137 251325 509149 251359
rect 509217 251325 509229 251359
rect 509137 251319 509229 251325
rect 509264 251233 509298 251397
rect 509346 251481 509380 251657
rect 509413 251553 509505 251559
rect 509413 251519 509425 251553
rect 509493 251519 509505 251553
rect 509413 251513 509505 251519
rect 509689 251553 509781 251559
rect 509689 251519 509701 251553
rect 509769 251519 509781 251553
rect 509689 251513 509781 251519
rect 509538 251481 509568 251493
rect 509346 251469 509403 251481
rect 509346 251409 509363 251469
rect 509397 251409 509403 251469
rect 509346 251397 509403 251409
rect 509515 251469 509568 251481
rect 509515 251409 509521 251469
rect 509555 251409 509568 251469
rect 509515 251397 509568 251409
rect 509346 251395 509380 251397
rect 509413 251359 509505 251365
rect 509413 251325 509425 251359
rect 509493 251325 509505 251359
rect 509413 251319 509505 251325
rect 509538 251233 509568 251397
rect 509626 251481 509656 251495
rect 509816 251481 509850 251657
rect 509626 251469 509679 251481
rect 509626 251409 509639 251469
rect 509673 251409 509679 251469
rect 509626 251397 509679 251409
rect 509791 251469 509850 251481
rect 509791 251409 509797 251469
rect 509831 251409 509850 251469
rect 509791 251397 509850 251409
rect 509902 251481 509936 251657
rect 509974 251595 510189 251605
rect 509974 251559 510104 251595
rect 509965 251553 510104 251559
rect 509965 251519 509977 251553
rect 510045 251535 510104 251553
rect 510164 251535 510189 251595
rect 510045 251525 510189 251535
rect 510241 251553 510333 251559
rect 510045 251519 510057 251525
rect 509965 251513 510057 251519
rect 510241 251519 510253 251553
rect 510321 251519 510333 251553
rect 510241 251513 510333 251519
rect 510086 251481 510116 251495
rect 509902 251469 509955 251481
rect 509902 251409 509915 251469
rect 509949 251409 509955 251469
rect 509902 251397 509955 251409
rect 510067 251469 510116 251481
rect 510067 251409 510073 251469
rect 510107 251409 510116 251469
rect 510067 251397 510116 251409
rect 509626 251233 509656 251397
rect 509902 251391 509936 251397
rect 509689 251359 509781 251365
rect 509689 251325 509701 251359
rect 509769 251325 509781 251359
rect 509965 251359 510057 251365
rect 509965 251340 509977 251359
rect 509689 251319 509781 251325
rect 509829 251335 509977 251340
rect 509829 251280 509839 251335
rect 509904 251325 509977 251335
rect 510045 251325 510057 251359
rect 509904 251319 510057 251325
rect 509904 251290 510044 251319
rect 509904 251280 509914 251290
rect 509829 251275 509914 251280
rect 510086 251233 510116 251397
rect 510178 251481 510208 251495
rect 510368 251481 510402 251657
rect 510178 251469 510231 251481
rect 510178 251409 510191 251469
rect 510225 251409 510231 251469
rect 510178 251397 510231 251409
rect 510343 251469 510402 251481
rect 510343 251409 510349 251469
rect 510383 251409 510402 251469
rect 510343 251399 510402 251409
rect 510454 251481 510488 251657
rect 510517 251553 510609 251559
rect 510517 251519 510529 251553
rect 510597 251519 510609 251553
rect 510517 251513 510609 251519
rect 510793 251553 510885 251559
rect 510793 251519 510805 251553
rect 510873 251519 510885 251553
rect 510793 251513 510885 251519
rect 510640 251481 510670 251495
rect 510454 251469 510507 251481
rect 510454 251409 510467 251469
rect 510501 251409 510507 251469
rect 510343 251397 510389 251399
rect 510454 251397 510507 251409
rect 510619 251469 510670 251481
rect 510619 251409 510625 251469
rect 510659 251409 510670 251469
rect 510619 251397 510670 251409
rect 510178 251233 510208 251397
rect 510454 251395 510488 251397
rect 510241 251359 510333 251365
rect 510241 251325 510253 251359
rect 510321 251325 510333 251359
rect 510241 251319 510333 251325
rect 510517 251359 510609 251365
rect 510517 251325 510529 251359
rect 510597 251325 510609 251359
rect 510517 251319 510609 251325
rect 510640 251233 510670 251397
rect 510732 251481 510762 251495
rect 510918 251481 510952 251657
rect 510732 251469 510783 251481
rect 510732 251409 510743 251469
rect 510777 251409 510783 251469
rect 510732 251397 510783 251409
rect 510895 251469 510952 251481
rect 510895 251409 510901 251469
rect 510935 251409 510952 251469
rect 510895 251397 510952 251409
rect 510732 251233 510762 251397
rect 510918 251395 510952 251397
rect 511006 251481 511040 251657
rect 511069 251553 511161 251559
rect 511069 251519 511081 251553
rect 511149 251519 511161 251553
rect 511069 251513 511161 251519
rect 511345 251553 511437 251559
rect 511345 251519 511357 251553
rect 511425 251519 511437 251553
rect 511345 251513 511437 251519
rect 511192 251481 511222 251495
rect 511006 251469 511059 251481
rect 511006 251409 511019 251469
rect 511053 251409 511059 251469
rect 511006 251397 511059 251409
rect 511171 251469 511222 251481
rect 511171 251409 511177 251469
rect 511211 251409 511222 251469
rect 511171 251397 511222 251409
rect 511006 251393 511040 251397
rect 510793 251359 510885 251365
rect 510793 251325 510805 251359
rect 510873 251325 510885 251359
rect 510793 251319 510885 251325
rect 511069 251359 511161 251365
rect 511069 251325 511081 251359
rect 511149 251325 511161 251359
rect 511069 251319 511161 251325
rect 511192 251233 511222 251397
rect 511278 251481 511308 251495
rect 511474 251481 511508 251657
rect 511278 251469 511335 251481
rect 511278 251409 511295 251469
rect 511329 251409 511335 251469
rect 511278 251397 511335 251409
rect 511447 251469 511508 251481
rect 511447 251409 511453 251469
rect 511487 251409 511508 251469
rect 511447 251397 511508 251409
rect 511278 251233 511308 251397
rect 511474 251389 511508 251397
rect 511556 251481 511590 251657
rect 511621 251553 511713 251559
rect 511621 251519 511633 251553
rect 511701 251519 511713 251553
rect 511621 251513 511713 251519
rect 511897 251553 511989 251559
rect 511897 251519 511909 251553
rect 511977 251519 511989 251553
rect 511897 251513 511989 251519
rect 511746 251481 511776 251495
rect 511556 251469 511611 251481
rect 511556 251409 511571 251469
rect 511605 251409 511611 251469
rect 511556 251397 511611 251409
rect 511723 251469 511776 251481
rect 511723 251409 511729 251469
rect 511763 251409 511776 251469
rect 511723 251397 511776 251409
rect 511556 251395 511590 251397
rect 511345 251359 511437 251365
rect 511345 251325 511357 251359
rect 511425 251325 511437 251359
rect 511345 251319 511437 251325
rect 511621 251359 511713 251365
rect 511621 251325 511633 251359
rect 511701 251325 511713 251359
rect 511621 251319 511713 251325
rect 511746 251233 511776 251397
rect 511834 251481 511864 251493
rect 512028 251481 512062 251657
rect 511834 251469 511887 251481
rect 511834 251409 511847 251469
rect 511881 251409 511887 251469
rect 511834 251397 511887 251409
rect 511999 251469 512062 251481
rect 511999 251409 512005 251469
rect 512039 251409 512062 251469
rect 511999 251397 512062 251409
rect 511834 251233 511864 251397
rect 512028 251393 512062 251397
rect 512106 251481 512140 251657
rect 512173 251553 512265 251559
rect 512173 251519 512185 251553
rect 512253 251519 512265 251553
rect 512173 251513 512265 251519
rect 512449 251553 512541 251559
rect 512449 251519 512461 251553
rect 512529 251519 512541 251553
rect 512449 251513 512541 251519
rect 512298 251481 512328 251497
rect 512106 251469 512163 251481
rect 512106 251409 512123 251469
rect 512157 251409 512163 251469
rect 512106 251397 512163 251409
rect 512275 251469 512328 251481
rect 512275 251409 512281 251469
rect 512315 251409 512328 251469
rect 512275 251397 512328 251409
rect 512106 251395 512140 251397
rect 511897 251359 511989 251365
rect 511897 251325 511909 251359
rect 511977 251325 511989 251359
rect 511897 251319 511989 251325
rect 512173 251359 512265 251365
rect 512173 251325 512185 251359
rect 512253 251325 512265 251359
rect 512173 251319 512265 251325
rect 512298 251233 512328 251397
rect 512386 251481 512416 251497
rect 512584 251481 512618 251657
rect 512386 251469 512439 251481
rect 512386 251409 512399 251469
rect 512433 251409 512439 251469
rect 512386 251397 512439 251409
rect 512551 251469 512618 251481
rect 512551 251409 512557 251469
rect 512591 251409 512618 251469
rect 512551 251397 512618 251409
rect 512386 251233 512416 251397
rect 512584 251385 512618 251397
rect 512658 251481 512692 251657
rect 512725 251553 512817 251559
rect 512725 251519 512737 251553
rect 512805 251519 512817 251553
rect 512725 251513 512817 251519
rect 513001 251553 513093 251559
rect 513001 251519 513013 251553
rect 513081 251519 513093 251553
rect 513001 251513 513093 251519
rect 512848 251481 512878 251499
rect 512658 251469 512715 251481
rect 512658 251409 512675 251469
rect 512709 251409 512715 251469
rect 512658 251397 512715 251409
rect 512827 251469 512878 251481
rect 512827 251409 512833 251469
rect 512867 251409 512878 251469
rect 512827 251397 512878 251409
rect 512658 251389 512692 251397
rect 512449 251359 512541 251365
rect 512449 251325 512461 251359
rect 512529 251325 512541 251359
rect 512449 251319 512541 251325
rect 512725 251359 512817 251365
rect 512725 251325 512737 251359
rect 512805 251325 512817 251359
rect 512725 251319 512817 251325
rect 512848 251233 512878 251397
rect 512936 251481 512966 251497
rect 513128 251481 513162 251657
rect 512936 251469 512991 251481
rect 512936 251409 512951 251469
rect 512985 251409 512991 251469
rect 512936 251397 512991 251409
rect 513103 251469 513162 251481
rect 513103 251409 513109 251469
rect 513143 251409 513162 251469
rect 513103 251397 513162 251409
rect 512936 251233 512966 251397
rect 513128 251385 513162 251397
rect 513208 251481 513242 251657
rect 513277 251553 513369 251559
rect 513277 251519 513289 251553
rect 513357 251519 513369 251553
rect 513277 251513 513369 251519
rect 513553 251553 513645 251559
rect 513553 251519 513565 251553
rect 513633 251519 513645 251553
rect 513553 251513 513645 251519
rect 513400 251481 513430 251497
rect 513208 251469 513267 251481
rect 513208 251409 513227 251469
rect 513261 251409 513267 251469
rect 513208 251397 513267 251409
rect 513379 251469 513430 251481
rect 513379 251409 513385 251469
rect 513419 251409 513430 251469
rect 513379 251397 513430 251409
rect 513208 251383 513242 251397
rect 513001 251359 513093 251365
rect 513001 251325 513013 251359
rect 513081 251325 513093 251359
rect 513001 251319 513093 251325
rect 513277 251359 513369 251365
rect 513277 251325 513289 251359
rect 513357 251325 513369 251359
rect 513277 251319 513369 251325
rect 513400 251233 513430 251397
rect 513488 251481 513518 251499
rect 513684 251481 513718 251657
rect 513488 251469 513543 251481
rect 513488 251409 513503 251469
rect 513537 251409 513543 251469
rect 513488 251397 513543 251409
rect 513655 251469 513718 251481
rect 513655 251409 513661 251469
rect 513695 251409 513718 251469
rect 513655 251397 513718 251409
rect 513488 251233 513518 251397
rect 513684 251385 513718 251397
rect 513758 251481 513792 251657
rect 513829 251553 513921 251559
rect 513829 251519 513841 251553
rect 513909 251519 513921 251553
rect 513829 251513 513921 251519
rect 514105 251553 514197 251559
rect 514105 251519 514117 251553
rect 514185 251519 514197 251553
rect 514105 251513 514197 251519
rect 513952 251481 513982 251497
rect 513758 251469 513819 251481
rect 513758 251409 513779 251469
rect 513813 251409 513819 251469
rect 513758 251397 513819 251409
rect 513931 251469 513982 251481
rect 513931 251409 513937 251469
rect 513971 251409 513982 251469
rect 513931 251397 513982 251409
rect 513758 251383 513792 251397
rect 513553 251359 513645 251365
rect 513553 251325 513565 251359
rect 513633 251325 513645 251359
rect 513553 251319 513645 251325
rect 513829 251359 513921 251365
rect 513829 251325 513841 251359
rect 513909 251325 513921 251359
rect 513829 251319 513921 251325
rect 513952 251233 513982 251397
rect 514042 251481 514072 251499
rect 514234 251481 514268 251657
rect 514042 251469 514095 251481
rect 514042 251409 514055 251469
rect 514089 251409 514095 251469
rect 514042 251397 514095 251409
rect 514207 251469 514268 251481
rect 514207 251409 514213 251469
rect 514247 251409 514268 251469
rect 514207 251397 514268 251409
rect 514042 251233 514072 251397
rect 514234 251387 514268 251397
rect 514310 251481 514344 251657
rect 514381 251553 514473 251559
rect 514381 251519 514393 251553
rect 514461 251519 514473 251553
rect 514381 251513 514473 251519
rect 514657 251553 514749 251559
rect 514657 251519 514669 251553
rect 514737 251519 514749 251553
rect 514657 251513 514749 251519
rect 514504 251481 514534 251497
rect 514310 251469 514371 251481
rect 514310 251409 514331 251469
rect 514365 251409 514371 251469
rect 514310 251397 514371 251409
rect 514483 251469 514534 251481
rect 514483 251409 514489 251469
rect 514523 251409 514534 251469
rect 514483 251397 514534 251409
rect 514310 251387 514344 251397
rect 514105 251359 514197 251365
rect 514105 251325 514117 251359
rect 514185 251325 514197 251359
rect 514105 251319 514197 251325
rect 514381 251359 514473 251365
rect 514381 251325 514393 251359
rect 514461 251325 514473 251359
rect 514381 251319 514473 251325
rect 514504 251233 514534 251397
rect 514594 251481 514624 251499
rect 514784 251481 514818 251657
rect 514594 251469 514647 251481
rect 514594 251409 514607 251469
rect 514641 251409 514647 251469
rect 514594 251397 514647 251409
rect 514759 251469 514818 251481
rect 514759 251409 514765 251469
rect 514799 251409 514818 251469
rect 514759 251397 514818 251409
rect 514594 251233 514624 251397
rect 514784 251391 514818 251397
rect 514866 251481 514900 251657
rect 514933 251553 515025 251559
rect 514933 251519 514945 251553
rect 515013 251519 515025 251553
rect 514933 251513 515025 251519
rect 515209 251553 515301 251559
rect 515209 251519 515221 251553
rect 515289 251519 515301 251553
rect 515209 251513 515301 251519
rect 515058 251481 515088 251503
rect 514866 251469 514923 251481
rect 514866 251409 514883 251469
rect 514917 251409 514923 251469
rect 514866 251397 514923 251409
rect 515035 251469 515088 251481
rect 515035 251409 515041 251469
rect 515075 251409 515088 251469
rect 515035 251397 515088 251409
rect 514866 251389 514900 251397
rect 514657 251359 514749 251365
rect 514657 251325 514669 251359
rect 514737 251325 514749 251359
rect 514657 251319 514749 251325
rect 514933 251359 515025 251365
rect 514933 251325 514945 251359
rect 515013 251325 515025 251359
rect 514933 251319 515025 251325
rect 515058 251233 515088 251397
rect 515148 251481 515178 251505
rect 515336 251481 515370 251657
rect 515148 251469 515199 251481
rect 515148 251409 515159 251469
rect 515193 251409 515199 251469
rect 515148 251397 515199 251409
rect 515311 251469 515370 251481
rect 515311 251409 515317 251469
rect 515351 251409 515370 251469
rect 515311 251397 515370 251409
rect 515414 251481 515448 251657
rect 515485 251553 515577 251559
rect 515485 251519 515497 251553
rect 515565 251519 515577 251553
rect 515485 251513 515577 251519
rect 515761 251553 515853 251559
rect 515761 251519 515773 251553
rect 515841 251519 515853 251553
rect 515761 251513 515853 251519
rect 515612 251481 515642 251505
rect 515414 251469 515475 251481
rect 515414 251409 515435 251469
rect 515469 251409 515475 251469
rect 515414 251397 515475 251409
rect 515587 251469 515642 251481
rect 515587 251409 515593 251469
rect 515627 251409 515642 251469
rect 515587 251397 515642 251409
rect 515148 251233 515178 251397
rect 515336 251395 515370 251397
rect 515209 251359 515301 251365
rect 515209 251325 515221 251359
rect 515289 251325 515301 251359
rect 515209 251319 515301 251325
rect 515485 251359 515577 251365
rect 515485 251325 515497 251359
rect 515565 251325 515577 251359
rect 515485 251319 515577 251325
rect 515612 251233 515642 251397
rect 515698 251481 515728 251509
rect 515886 251481 515920 251657
rect 515698 251469 515751 251481
rect 515698 251409 515711 251469
rect 515745 251409 515751 251469
rect 515698 251397 515751 251409
rect 515863 251469 515920 251481
rect 515863 251409 515869 251469
rect 515903 251409 515920 251469
rect 515863 251397 515920 251409
rect 515698 251233 515728 251397
rect 515886 251393 515920 251397
rect 515970 251481 516004 251657
rect 516037 251553 516129 251559
rect 516037 251519 516049 251553
rect 516117 251519 516129 251553
rect 516037 251513 516129 251519
rect 516313 251553 516405 251559
rect 516313 251519 516325 251553
rect 516393 251519 516405 251553
rect 516313 251513 516405 251519
rect 516158 251481 516188 251495
rect 515970 251469 516027 251481
rect 515970 251409 515987 251469
rect 516021 251409 516027 251469
rect 515970 251397 516027 251409
rect 516139 251469 516188 251481
rect 516139 251409 516145 251469
rect 516179 251409 516188 251469
rect 516139 251397 516188 251409
rect 515970 251391 516004 251397
rect 515761 251359 515853 251365
rect 515761 251325 515773 251359
rect 515841 251325 515853 251359
rect 515761 251319 515853 251325
rect 516037 251359 516129 251365
rect 516037 251325 516049 251359
rect 516117 251325 516129 251359
rect 516037 251319 516129 251325
rect 516158 251233 516188 251397
rect 516250 251481 516280 251493
rect 516438 251481 516472 251657
rect 516250 251469 516303 251481
rect 516250 251409 516263 251469
rect 516297 251409 516303 251469
rect 516250 251397 516303 251409
rect 516415 251469 516472 251481
rect 516415 251409 516421 251469
rect 516455 251409 516472 251469
rect 516415 251397 516472 251409
rect 516250 251233 516280 251397
rect 516438 251393 516472 251397
rect 516522 251481 516556 251657
rect 516589 251553 516681 251559
rect 516589 251519 516601 251553
rect 516669 251519 516681 251553
rect 516589 251513 516681 251519
rect 516865 251553 516957 251559
rect 516865 251519 516877 251553
rect 516945 251519 516957 251553
rect 516865 251513 516957 251519
rect 516714 251481 516744 251495
rect 516522 251469 516579 251481
rect 516522 251409 516539 251469
rect 516573 251409 516579 251469
rect 516522 251397 516579 251409
rect 516691 251469 516744 251481
rect 516691 251409 516697 251469
rect 516731 251409 516744 251469
rect 516691 251397 516744 251409
rect 516522 251395 516556 251397
rect 516313 251359 516405 251365
rect 516313 251325 516325 251359
rect 516393 251325 516405 251359
rect 516313 251319 516405 251325
rect 516589 251359 516681 251365
rect 516589 251325 516601 251359
rect 516669 251325 516681 251359
rect 516589 251319 516681 251325
rect 516714 251233 516744 251397
rect 516798 251481 516828 251495
rect 516992 251481 517026 251657
rect 516798 251469 516855 251481
rect 516798 251409 516815 251469
rect 516849 251409 516855 251469
rect 516798 251397 516855 251409
rect 516967 251469 517026 251481
rect 516967 251409 516973 251469
rect 517007 251409 517026 251469
rect 516967 251399 517026 251409
rect 517070 251481 517104 251657
rect 517141 251553 517233 251559
rect 517141 251519 517153 251553
rect 517221 251519 517233 251553
rect 517141 251513 517233 251519
rect 517264 251481 517294 251495
rect 517070 251469 517131 251481
rect 517070 251409 517091 251469
rect 517125 251409 517131 251469
rect 516967 251397 517013 251399
rect 517070 251397 517131 251409
rect 517243 251469 517294 251481
rect 517243 251409 517249 251469
rect 517283 251409 517294 251469
rect 517243 251397 517294 251409
rect 517384 251405 517418 251657
rect 516798 251233 516828 251397
rect 516865 251359 516957 251365
rect 516865 251325 516877 251359
rect 516945 251325 516957 251359
rect 516865 251319 516957 251325
rect 517141 251359 517233 251365
rect 517141 251325 517153 251359
rect 517221 251325 517233 251359
rect 517141 251319 517233 251325
rect 517264 251233 517294 251397
rect 503127 251191 517296 251233
rect 517254 251189 517296 251191
rect 507306 251085 507446 251097
rect 507306 251029 507346 251085
rect 507424 251029 507446 251085
rect 507306 250415 507446 251029
rect 518318 250600 519188 251657
rect 501258 248634 502348 248640
rect 503138 250215 507492 250415
rect 503138 245815 503338 250215
rect 518318 249724 519188 249730
rect 322310 239406 322640 240230
rect 323366 239406 323762 240230
rect 322310 238812 323762 239406
rect 412310 240230 413762 245815
rect 412310 239406 412640 240230
rect 413366 239406 413762 240230
rect 412310 238812 413762 239406
rect 502310 240230 503762 245815
rect 502310 239406 502640 240230
rect 503366 239406 503762 240230
rect 502310 238812 503762 239406
rect 57138 149300 58098 149460
rect 57138 148700 57298 149300
rect 57898 148700 58098 149300
rect 57138 147780 58098 148700
rect 60858 149300 61818 149460
rect 60858 148700 61018 149300
rect 61618 148700 61818 149300
rect 60858 147780 61818 148700
rect 57138 147180 61818 147780
rect 147138 149300 148098 149460
rect 147138 148700 147298 149300
rect 147898 148700 148098 149300
rect 147138 147780 148098 148700
rect 150858 149300 151818 149460
rect 150858 148700 151018 149300
rect 151618 148700 151818 149300
rect 150858 147780 151818 148700
rect 147138 147180 151818 147780
rect 237138 149300 238098 149460
rect 237138 148700 237298 149300
rect 237898 148700 238098 149300
rect 237138 147780 238098 148700
rect 240858 149300 241818 149460
rect 240858 148700 241018 149300
rect 241618 148700 241818 149300
rect 240858 147780 241818 148700
rect 237138 147180 241818 147780
rect 327138 149300 328098 149460
rect 327138 148700 327298 149300
rect 327898 148700 328098 149300
rect 327138 147780 328098 148700
rect 330858 149300 331818 149460
rect 330858 148700 331018 149300
rect 331618 148700 331818 149300
rect 330858 147780 331818 148700
rect 327138 147180 331818 147780
rect 417138 149300 418098 149460
rect 417138 148700 417298 149300
rect 417898 148700 418098 149300
rect 417138 147780 418098 148700
rect 420858 149300 421818 149460
rect 420858 148700 421018 149300
rect 421618 148700 421818 149300
rect 420858 147780 421818 148700
rect 417138 147180 421818 147780
rect 507138 149300 508098 149460
rect 507138 148700 507298 149300
rect 507898 148700 508098 149300
rect 507138 147780 508098 148700
rect 510858 149300 511818 149460
rect 510858 148700 511018 149300
rect 511618 148700 511818 149300
rect 510858 147780 511818 148700
rect 507138 147180 511818 147780
rect 59258 146320 59498 147180
rect 59338 146033 59378 146320
rect 149458 146300 149658 147180
rect 239238 146760 239440 147180
rect 239238 146578 239438 146760
rect 59327 146027 59385 146033
rect 58118 145980 58558 146000
rect 59327 145993 59339 146027
rect 59373 145993 59385 146027
rect 59327 145987 59385 145993
rect 58118 145960 58918 145980
rect 58118 145800 58178 145960
rect 58338 145900 58918 145960
rect 60078 145960 60558 145980
rect 59289 145934 59335 145946
rect 59289 145900 59295 145934
rect 58338 145840 59295 145900
rect 58338 145800 58918 145840
rect 58118 145760 58918 145800
rect 59289 145758 59295 145840
rect 59329 145758 59335 145934
rect 59289 145746 59335 145758
rect 59377 145934 59423 145946
rect 59377 145758 59383 145934
rect 59417 145900 59423 145934
rect 60078 145900 60378 145960
rect 59417 145840 60378 145900
rect 59417 145758 59423 145840
rect 60078 145800 60378 145840
rect 60538 145800 60558 145960
rect 60078 145780 60558 145800
rect 148118 145960 148858 146000
rect 148118 145800 148178 145960
rect 148338 145800 148858 145960
rect 148118 145760 148858 145800
rect 59377 145746 59423 145758
rect 59327 145699 59385 145705
rect 59327 145665 59339 145699
rect 59373 145665 59385 145699
rect 59327 145659 59385 145665
rect 59338 145380 59378 145659
rect 148658 145540 148858 145760
rect 149518 145623 149638 146300
rect 239298 146056 239438 146578
rect 329258 146320 329498 147180
rect 239298 146038 239356 146056
rect 239340 146022 239356 146038
rect 239390 146038 239438 146056
rect 239390 146022 239402 146038
rect 329338 146033 329378 146320
rect 419458 146300 419658 147180
rect 509238 146760 509440 147180
rect 509238 146578 509438 146760
rect 239340 146020 239402 146022
rect 239344 146016 239402 146020
rect 329327 146027 329385 146033
rect 149518 145589 149537 145623
rect 149605 145589 149638 145623
rect 149518 145580 149638 145589
rect 150358 145960 150558 145980
rect 150358 145800 150378 145960
rect 150538 145800 150558 145960
rect 149469 145540 149515 145542
rect 148658 145530 149515 145540
rect 59278 144240 59498 145380
rect 148658 145354 149475 145530
rect 149509 145354 149515 145530
rect 148658 145342 149515 145354
rect 149627 145540 149673 145542
rect 150358 145540 150558 145800
rect 238118 145960 238918 146000
rect 238118 145800 238178 145960
rect 238338 145940 238918 145960
rect 239306 145972 239352 145984
rect 239306 145940 239312 145972
rect 238338 145820 239312 145940
rect 238338 145800 238918 145820
rect 238118 145760 238918 145800
rect 239306 145796 239312 145820
rect 239346 145796 239352 145972
rect 239306 145784 239352 145796
rect 239394 145972 239440 145984
rect 328118 145980 328558 146000
rect 329327 145993 329339 146027
rect 329373 145993 329385 146027
rect 329327 145987 329385 145993
rect 239394 145796 239400 145972
rect 239434 145940 239440 145972
rect 240358 145960 240558 145980
rect 240358 145940 240378 145960
rect 239434 145820 240378 145940
rect 239434 145796 239440 145820
rect 239394 145784 239440 145796
rect 240358 145800 240378 145820
rect 240538 145800 240558 145960
rect 240358 145780 240558 145800
rect 328118 145960 328918 145980
rect 328118 145800 328178 145960
rect 328338 145900 328918 145960
rect 330078 145960 330558 145980
rect 329289 145934 329335 145946
rect 329289 145900 329295 145934
rect 328338 145840 329295 145900
rect 328338 145800 328918 145840
rect 328118 145760 328918 145800
rect 329289 145758 329295 145840
rect 329329 145758 329335 145934
rect 239344 145746 239402 145752
rect 329289 145746 329335 145758
rect 329377 145934 329423 145946
rect 329377 145758 329383 145934
rect 329417 145900 329423 145934
rect 330078 145900 330378 145960
rect 329417 145840 330378 145900
rect 329417 145758 329423 145840
rect 330078 145800 330378 145840
rect 330538 145800 330558 145960
rect 330078 145780 330558 145800
rect 418118 145960 418858 146000
rect 418118 145800 418178 145960
rect 418338 145800 418858 145960
rect 418118 145760 418858 145800
rect 329377 145746 329423 145758
rect 239344 145740 239356 145746
rect 149627 145530 150558 145540
rect 149627 145354 149633 145530
rect 149667 145354 150558 145530
rect 149627 145342 150558 145354
rect 148658 145340 149498 145342
rect 149638 145340 150558 145342
rect 239298 145712 239356 145740
rect 239390 145740 239402 145746
rect 239390 145712 239438 145740
rect 149525 145300 149617 145301
rect 149518 145295 149618 145300
rect 149518 145261 149537 145295
rect 149605 145261 149618 145295
rect 149518 144840 149618 145261
rect 239298 145200 239438 145712
rect 329327 145699 329385 145705
rect 329327 145665 329339 145699
rect 329373 145665 329385 145699
rect 329327 145659 329385 145665
rect 329338 145380 329378 145659
rect 418658 145540 418858 145760
rect 419518 145623 419638 146300
rect 509298 146056 509438 146578
rect 509298 146038 509356 146056
rect 509340 146022 509356 146038
rect 509390 146038 509438 146056
rect 509390 146022 509402 146038
rect 509340 146020 509402 146022
rect 509344 146016 509402 146020
rect 419518 145589 419537 145623
rect 419605 145589 419638 145623
rect 419518 145580 419638 145589
rect 420358 145960 420558 145980
rect 420358 145800 420378 145960
rect 420538 145800 420558 145960
rect 419469 145540 419515 145542
rect 418658 145530 419515 145540
rect 149458 144240 149658 144840
rect 239238 144240 239438 145200
rect 329278 144240 329498 145380
rect 418658 145354 419475 145530
rect 419509 145354 419515 145530
rect 418658 145342 419515 145354
rect 419627 145540 419673 145542
rect 420358 145540 420558 145800
rect 508118 145960 508918 146000
rect 508118 145800 508178 145960
rect 508338 145940 508918 145960
rect 509306 145972 509352 145984
rect 509306 145940 509312 145972
rect 508338 145820 509312 145940
rect 508338 145800 508918 145820
rect 508118 145760 508918 145800
rect 509306 145796 509312 145820
rect 509346 145796 509352 145972
rect 509306 145784 509352 145796
rect 509394 145972 509440 145984
rect 509394 145796 509400 145972
rect 509434 145940 509440 145972
rect 510358 145960 510558 145980
rect 510358 145940 510378 145960
rect 509434 145820 510378 145940
rect 509434 145796 509440 145820
rect 509394 145784 509440 145796
rect 510358 145800 510378 145820
rect 510538 145800 510558 145960
rect 510358 145780 510558 145800
rect 509344 145746 509402 145752
rect 509344 145740 509356 145746
rect 419627 145530 420558 145540
rect 419627 145354 419633 145530
rect 419667 145354 420558 145530
rect 419627 145342 420558 145354
rect 418658 145340 419498 145342
rect 419638 145340 420558 145342
rect 509298 145712 509356 145740
rect 509390 145740 509402 145746
rect 509390 145712 509438 145740
rect 419525 145300 419617 145301
rect 419518 145295 419618 145300
rect 419518 145261 419537 145295
rect 419605 145261 419618 145295
rect 419518 144840 419618 145261
rect 509298 145200 509438 145712
rect 419458 144240 419658 144840
rect 509238 144240 509438 145200
rect 57078 143640 61758 144240
rect 57078 142720 58038 143640
rect 57078 142120 57238 142720
rect 57838 142120 58038 142720
rect 57078 141960 58038 142120
rect 60798 142720 61758 143640
rect 60798 142120 60958 142720
rect 61558 142120 61758 142720
rect 60798 141960 61758 142120
rect 147078 143640 151758 144240
rect 147078 142720 148038 143640
rect 147078 142120 147238 142720
rect 147838 142120 148038 142720
rect 147078 141960 148038 142120
rect 150798 142720 151758 143640
rect 150798 142120 150958 142720
rect 151558 142120 151758 142720
rect 150798 141960 151758 142120
rect 237078 143640 241758 144240
rect 237078 142720 238038 143640
rect 237078 142120 237238 142720
rect 237838 142120 238038 142720
rect 237078 141960 238038 142120
rect 240798 142720 241758 143640
rect 240798 142120 240958 142720
rect 241558 142120 241758 142720
rect 240798 141960 241758 142120
rect 327078 143640 331758 144240
rect 327078 142720 328038 143640
rect 327078 142120 327238 142720
rect 327838 142120 328038 142720
rect 327078 141960 328038 142120
rect 330798 142720 331758 143640
rect 330798 142120 330958 142720
rect 331558 142120 331758 142720
rect 330798 141960 331758 142120
rect 417078 143640 421758 144240
rect 417078 142720 418038 143640
rect 417078 142120 417238 142720
rect 417838 142120 418038 142720
rect 417078 141960 418038 142120
rect 420798 142720 421758 143640
rect 420798 142120 420958 142720
rect 421558 142120 421758 142720
rect 420798 141960 421758 142120
rect 507078 143640 511758 144240
rect 507078 142720 508038 143640
rect 507078 142120 507238 142720
rect 507838 142120 508038 142720
rect 507078 141960 508038 142120
rect 510798 142720 511758 143640
rect 510798 142120 510958 142720
rect 511558 142120 511758 142720
rect 510798 141960 511758 142120
rect 57138 59300 58098 59460
rect 57138 58700 57298 59300
rect 57898 58700 58098 59300
rect 57138 57780 58098 58700
rect 60858 59300 61818 59460
rect 60858 58700 61018 59300
rect 61618 58700 61818 59300
rect 60858 57780 61818 58700
rect 57138 57180 61818 57780
rect 147138 59300 148098 59460
rect 147138 58700 147298 59300
rect 147898 58700 148098 59300
rect 147138 57780 148098 58700
rect 150858 59300 151818 59460
rect 150858 58700 151018 59300
rect 151618 58700 151818 59300
rect 149198 57780 149498 57790
rect 150858 57780 151818 58700
rect 147138 57190 151818 57780
rect 147138 57180 149238 57190
rect 149498 57180 151818 57190
rect 237138 59300 238098 59460
rect 237138 58700 237298 59300
rect 237898 58700 238098 59300
rect 237138 57780 238098 58700
rect 240858 59300 241818 59460
rect 240858 58700 241018 59300
rect 241618 58700 241818 59300
rect 240858 57780 241818 58700
rect 237138 57180 241818 57780
rect 327138 59300 328098 59460
rect 327138 58700 327298 59300
rect 327898 58700 328098 59300
rect 327138 57780 328098 58700
rect 330858 59300 331818 59460
rect 330858 58700 331018 59300
rect 331618 58700 331818 59300
rect 330858 57780 331818 58700
rect 327138 57180 331818 57780
rect 417138 59300 418098 59460
rect 417138 58700 417298 59300
rect 417898 58700 418098 59300
rect 417138 57780 418098 58700
rect 420858 59300 421818 59460
rect 420858 58700 421018 59300
rect 421618 58700 421818 59300
rect 419198 57780 419498 57790
rect 420858 57780 421818 58700
rect 417138 57190 421818 57780
rect 417138 57180 419238 57190
rect 419498 57180 421818 57190
rect 507138 59300 508098 59460
rect 507138 58700 507298 59300
rect 507898 58700 508098 59300
rect 507138 57780 508098 58700
rect 510858 59300 511818 59460
rect 510858 58700 511018 59300
rect 511618 58700 511818 59300
rect 510858 57780 511818 58700
rect 507138 57180 511818 57780
rect 59238 56760 59440 57180
rect 59238 56578 59438 56760
rect 149548 56640 149748 57180
rect 59298 56056 59438 56578
rect 59298 56038 59356 56056
rect 59340 56022 59356 56038
rect 59390 56038 59438 56056
rect 149598 56061 149698 56640
rect 239558 56520 239778 57180
rect 329238 56760 329440 57180
rect 329238 56578 329438 56760
rect 419548 56640 419748 57180
rect 149598 56055 149707 56061
rect 149598 56040 149627 56055
rect 59390 56022 59402 56038
rect 59340 56020 59402 56022
rect 59344 56016 59402 56020
rect 149615 56021 149627 56040
rect 149695 56021 149707 56055
rect 149615 56015 149707 56021
rect 58118 55960 58918 56000
rect 58118 55800 58178 55960
rect 58338 55940 58918 55960
rect 59306 55972 59352 55984
rect 59306 55940 59312 55972
rect 58338 55820 59312 55940
rect 58338 55800 58918 55820
rect 58118 55760 58918 55800
rect 59306 55796 59312 55820
rect 59346 55796 59352 55972
rect 59306 55784 59352 55796
rect 59394 55972 59440 55984
rect 59394 55796 59400 55972
rect 59434 55940 59440 55972
rect 60358 55960 60558 55980
rect 60358 55940 60378 55960
rect 59434 55820 60378 55940
rect 59434 55796 59440 55820
rect 59394 55784 59440 55796
rect 60358 55800 60378 55820
rect 60538 55800 60558 55960
rect 60358 55780 60558 55800
rect 148118 55960 148918 56000
rect 148118 55800 148178 55960
rect 148338 55940 148918 55960
rect 149559 55971 149605 55983
rect 149559 55940 149565 55971
rect 148338 55840 149565 55940
rect 148338 55800 148918 55840
rect 148118 55760 148918 55800
rect 149559 55795 149565 55840
rect 149599 55795 149605 55971
rect 149559 55783 149605 55795
rect 149717 55971 149763 55983
rect 149717 55795 149723 55971
rect 149757 55940 149763 55971
rect 150348 55960 150548 55990
rect 150348 55940 150378 55960
rect 149757 55840 150378 55940
rect 149757 55795 149763 55840
rect 149717 55783 149763 55795
rect 150348 55800 150378 55840
rect 150538 55800 150548 55960
rect 150348 55790 150548 55800
rect 238118 55960 238858 56000
rect 238118 55800 238178 55960
rect 238338 55800 238858 55960
rect 238118 55760 238858 55800
rect 59344 55746 59402 55752
rect 59344 55740 59356 55746
rect 59298 55712 59356 55740
rect 59390 55740 59402 55746
rect 149615 55745 149707 55751
rect 149615 55740 149627 55745
rect 59390 55712 59438 55740
rect 59298 55200 59438 55712
rect 149598 55711 149627 55740
rect 149695 55711 149707 55745
rect 149598 55705 149707 55711
rect 149598 55290 149698 55705
rect 238658 55660 238858 55760
rect 239618 55765 239718 56520
rect 329298 56056 329438 56578
rect 329298 56038 329356 56056
rect 329340 56022 329356 56038
rect 329390 56038 329438 56056
rect 419598 56061 419698 56640
rect 509558 56520 509778 57180
rect 419598 56055 419707 56061
rect 419598 56040 419627 56055
rect 329390 56022 329402 56038
rect 329340 56020 329402 56022
rect 329344 56016 329402 56020
rect 419615 56021 419627 56040
rect 419695 56021 419707 56055
rect 419615 56015 419707 56021
rect 239618 55740 239637 55765
rect 239625 55731 239637 55740
rect 239705 55740 239718 55765
rect 240358 55960 240558 55980
rect 240358 55800 240378 55960
rect 240538 55800 240558 55960
rect 239705 55731 239717 55740
rect 239625 55725 239717 55731
rect 239569 55681 239615 55693
rect 239569 55660 239575 55681
rect 238658 55560 239575 55660
rect 238658 55500 238858 55560
rect 239569 55505 239575 55560
rect 239609 55505 239615 55681
rect 239569 55493 239615 55505
rect 239727 55681 239773 55693
rect 239727 55505 239733 55681
rect 239767 55660 239773 55681
rect 240358 55660 240558 55800
rect 328118 55960 328918 56000
rect 328118 55800 328178 55960
rect 328338 55940 328918 55960
rect 329306 55972 329352 55984
rect 329306 55940 329312 55972
rect 328338 55820 329312 55940
rect 328338 55800 328918 55820
rect 328118 55760 328918 55800
rect 329306 55796 329312 55820
rect 329346 55796 329352 55972
rect 329306 55784 329352 55796
rect 329394 55972 329440 55984
rect 329394 55796 329400 55972
rect 329434 55940 329440 55972
rect 330358 55960 330558 55980
rect 330358 55940 330378 55960
rect 329434 55820 330378 55940
rect 329434 55796 329440 55820
rect 329394 55784 329440 55796
rect 330358 55800 330378 55820
rect 330538 55800 330558 55960
rect 330358 55780 330558 55800
rect 418118 55960 418918 56000
rect 418118 55800 418178 55960
rect 418338 55940 418918 55960
rect 419559 55971 419605 55983
rect 419559 55940 419565 55971
rect 418338 55840 419565 55940
rect 418338 55800 418918 55840
rect 418118 55760 418918 55800
rect 419559 55795 419565 55840
rect 419599 55795 419605 55971
rect 419559 55783 419605 55795
rect 419717 55971 419763 55983
rect 419717 55795 419723 55971
rect 419757 55940 419763 55971
rect 420348 55960 420548 55990
rect 420348 55940 420378 55960
rect 419757 55840 420378 55940
rect 419757 55795 419763 55840
rect 419717 55783 419763 55795
rect 420348 55800 420378 55840
rect 420538 55800 420548 55960
rect 420348 55790 420548 55800
rect 508118 55960 508858 56000
rect 508118 55800 508178 55960
rect 508338 55800 508858 55960
rect 508118 55760 508858 55800
rect 329344 55746 329402 55752
rect 329344 55740 329356 55746
rect 239767 55560 240558 55660
rect 239767 55505 239773 55560
rect 239727 55493 239773 55505
rect 240358 55500 240558 55560
rect 329298 55712 329356 55740
rect 329390 55740 329402 55746
rect 419615 55745 419707 55751
rect 419615 55740 419627 55745
rect 329390 55712 329438 55740
rect 239625 55460 239717 55461
rect 239618 55455 239717 55460
rect 239618 55421 239637 55455
rect 239705 55421 239717 55455
rect 239618 55415 239717 55421
rect 59238 54240 59438 55200
rect 149548 54240 149748 55290
rect 239618 54900 239698 55415
rect 329298 55200 329438 55712
rect 419598 55711 419627 55740
rect 419695 55711 419707 55745
rect 419598 55705 419707 55711
rect 419598 55290 419698 55705
rect 508658 55660 508858 55760
rect 509618 55765 509718 56520
rect 509618 55740 509637 55765
rect 509625 55731 509637 55740
rect 509705 55740 509718 55765
rect 510358 55960 510558 55980
rect 510358 55800 510378 55960
rect 510538 55800 510558 55960
rect 509705 55731 509717 55740
rect 509625 55725 509717 55731
rect 509569 55681 509615 55693
rect 509569 55660 509575 55681
rect 508658 55560 509575 55660
rect 508658 55500 508858 55560
rect 509569 55505 509575 55560
rect 509609 55505 509615 55681
rect 509569 55493 509615 55505
rect 509727 55681 509773 55693
rect 509727 55505 509733 55681
rect 509767 55660 509773 55681
rect 510358 55660 510558 55800
rect 509767 55560 510558 55660
rect 509767 55505 509773 55560
rect 509727 55493 509773 55505
rect 510358 55500 510558 55560
rect 509625 55460 509717 55461
rect 509618 55455 509717 55460
rect 509618 55421 509637 55455
rect 509705 55421 509717 55455
rect 509618 55415 509717 55421
rect 239558 54240 239758 54900
rect 329238 54240 329438 55200
rect 419548 54240 419748 55290
rect 509618 54900 509698 55415
rect 509558 54240 509758 54900
rect 57078 53640 61758 54240
rect 57078 52720 58038 53640
rect 57078 52120 57238 52720
rect 57838 52120 58038 52720
rect 57078 51960 58038 52120
rect 60798 52720 61758 53640
rect 60798 52120 60958 52720
rect 61558 52120 61758 52720
rect 60798 51960 61758 52120
rect 147078 53640 151758 54240
rect 147078 52720 148038 53640
rect 147078 52120 147238 52720
rect 147838 52120 148038 52720
rect 147078 51960 148038 52120
rect 150798 52720 151758 53640
rect 150798 52120 150958 52720
rect 151558 52120 151758 52720
rect 150798 51960 151758 52120
rect 237078 53640 241758 54240
rect 237078 52720 238038 53640
rect 237078 52120 237238 52720
rect 237838 52120 238038 52720
rect 237078 51960 238038 52120
rect 240798 52720 241758 53640
rect 240798 52120 240958 52720
rect 241558 52120 241758 52720
rect 240798 51960 241758 52120
rect 327078 53640 331758 54240
rect 327078 52720 328038 53640
rect 327078 52120 327238 52720
rect 327838 52120 328038 52720
rect 327078 51960 328038 52120
rect 330798 52720 331758 53640
rect 330798 52120 330958 52720
rect 331558 52120 331758 52720
rect 330798 51960 331758 52120
rect 417078 53640 421758 54240
rect 417078 52720 418038 53640
rect 417078 52120 417238 52720
rect 417838 52120 418038 52720
rect 417078 51960 418038 52120
rect 420798 52720 421758 53640
rect 420798 52120 420958 52720
rect 421558 52120 421758 52720
rect 420798 51960 421758 52120
rect 507078 53640 511758 54240
rect 507078 52720 508038 53640
rect 507078 52120 507238 52720
rect 507838 52120 508038 52720
rect 507078 51960 508038 52120
rect 510798 52720 511758 53640
rect 510798 52120 510958 52720
rect 511558 52120 511758 52720
rect 510798 51960 511758 52120
<< via1 >>
rect 327100 660624 327700 661224
rect 330820 660624 331420 661224
rect 57298 658700 57898 659300
rect 61018 658700 61618 659300
rect 147298 658700 147898 659300
rect 151018 658700 151618 659300
rect 237298 658700 237898 659300
rect 241018 658700 241618 659300
rect 417100 660624 417700 661224
rect 420820 660624 421420 661224
rect 507100 660624 507700 661224
rect 510820 660624 511420 661224
rect 327980 657724 328140 657884
rect 330180 657724 330340 657884
rect 417980 657724 418140 657884
rect 420180 657724 420340 657884
rect 507980 657724 508140 657884
rect 510180 657724 510340 657884
rect 58178 655800 58338 655960
rect 60378 655800 60538 655960
rect 148178 655800 148338 655960
rect 150378 655800 150538 655960
rect 238178 655800 238338 655960
rect 240378 655800 240538 655960
rect 57238 652120 57838 652720
rect 60958 652120 61558 652720
rect 147238 652120 147838 652720
rect 150958 652120 151558 652720
rect 327040 654044 327640 654644
rect 330760 654044 331360 654644
rect 417040 654044 417640 654644
rect 420760 654044 421360 654644
rect 507040 654044 507640 654644
rect 510760 654044 511360 654644
rect 237238 652120 237838 652720
rect 240958 652120 241558 652720
rect 417100 585624 417700 586224
rect 420820 585624 421420 586224
rect 57298 583700 57898 584300
rect 61018 583700 61618 584300
rect 147298 583700 147898 584300
rect 151018 583700 151618 584300
rect 237298 583700 237898 584300
rect 241018 583700 241618 584300
rect 327298 583700 327898 584300
rect 331018 583700 331618 584300
rect 507100 585624 507700 586224
rect 510820 585624 511420 586224
rect 417980 582724 418140 582884
rect 420180 582724 420340 582884
rect 507980 582724 508140 582884
rect 510180 582724 510340 582884
rect 58178 580800 58338 580960
rect 60378 580800 60538 580960
rect 148178 580800 148338 580960
rect 150378 580800 150538 580960
rect 238178 580800 238338 580960
rect 240378 580800 240538 580960
rect 328178 580800 328338 580960
rect 330378 580800 330538 580960
rect 57238 577120 57838 577720
rect 60958 577120 61558 577720
rect 147238 577120 147838 577720
rect 150958 577120 151558 577720
rect 237238 577120 237838 577720
rect 240958 577120 241558 577720
rect 417040 579044 417640 579644
rect 420760 579044 421360 579644
rect 507040 579044 507640 579644
rect 510760 579044 511360 579644
rect 327238 577120 327838 577720
rect 330958 577120 331558 577720
rect 64790 503970 65516 504794
rect 57298 494800 57898 495400
rect 61018 494800 61618 495400
rect 154790 503970 155516 504794
rect 244790 503970 245516 504794
rect 334790 503970 335516 504794
rect 424790 503970 425516 504794
rect 417298 494800 417898 495400
rect 421018 494800 421618 495400
rect 514790 503970 515516 504794
rect 323908 493378 324016 493502
rect 60008 492328 60080 492392
rect 57996 491684 58146 491786
rect 60008 491843 60076 491872
rect 60008 491816 60075 491843
rect 60075 491816 60076 491843
rect 60008 491615 60075 491642
rect 60075 491615 60076 491642
rect 60008 491586 60076 491615
rect 62696 491638 62844 491786
rect 230433 491842 231381 492790
rect 507298 494800 507898 495400
rect 511018 494800 511618 495400
rect 321793 492028 322119 492354
rect 60012 491206 60084 491270
rect 57238 488220 57838 488820
rect 60958 488220 61558 488820
rect 150104 491535 150164 491595
rect 149839 491280 149904 491335
rect 323896 491500 323964 491556
rect 418178 491900 418338 492060
rect 510008 492328 510080 492392
rect 338860 491364 339000 491610
rect 419441 491784 419535 491844
rect 420378 491900 420538 492060
rect 141258 488640 142348 489730
rect 158318 489730 159188 490600
rect 239461 490939 239521 490999
rect 239196 490684 239261 490739
rect 247591 488633 249092 490134
rect 419445 491515 419531 491542
rect 419445 491484 419454 491515
rect 419454 491484 419522 491515
rect 419522 491484 419531 491515
rect 419445 491287 419454 491318
rect 419454 491287 419522 491318
rect 419522 491287 419531 491318
rect 419445 491260 419531 491287
rect 507996 491684 508146 491786
rect 510008 491843 510076 491872
rect 510008 491816 510075 491843
rect 510075 491816 510076 491843
rect 510008 491615 510075 491642
rect 510075 491615 510076 491642
rect 510008 491586 510076 491615
rect 512696 491638 512844 491786
rect 510012 491206 510084 491270
rect 419439 490930 419533 490990
rect 52640 479406 53366 480230
rect 142640 479406 143366 480230
rect 232640 479406 233366 480230
rect 322640 479406 323366 480230
rect 417238 488220 417838 488820
rect 420958 488220 421558 488820
rect 412640 479406 413366 480230
rect 507238 488220 507838 488820
rect 510958 488220 511558 488820
rect 502640 479406 503366 480230
rect 64790 383970 65516 384794
rect 154790 383970 155516 384794
rect 244790 383970 245516 384794
rect 334790 383970 335516 384794
rect 424790 383970 425516 384794
rect 417298 374800 417898 375400
rect 421018 374800 421618 375400
rect 514790 383970 515516 384794
rect 323908 373378 324016 373502
rect 60104 371535 60164 371595
rect 59839 371280 59904 371335
rect 51258 368640 52348 369730
rect 68318 369730 69188 370600
rect 230433 371842 231381 372790
rect 507298 374800 507898 375400
rect 511018 374800 511618 375400
rect 321793 372028 322119 372354
rect 150104 371535 150164 371595
rect 149839 371280 149904 371335
rect 323896 371500 323964 371556
rect 420008 372328 420080 372392
rect 417996 371684 418146 371786
rect 338860 371364 339000 371610
rect 420008 371843 420076 371872
rect 420008 371816 420075 371843
rect 420075 371816 420076 371843
rect 420008 371615 420075 371642
rect 420075 371615 420076 371642
rect 420008 371586 420076 371615
rect 508178 371900 508338 372060
rect 422696 371638 422844 371786
rect 509441 371784 509535 371844
rect 510378 371900 510538 372060
rect 420012 371206 420084 371270
rect 141258 368640 142348 369730
rect 158318 369730 159188 370600
rect 239461 370939 239521 370999
rect 239196 370684 239261 370739
rect 247591 368633 249092 370134
rect 509445 371515 509531 371542
rect 509445 371484 509454 371515
rect 509454 371484 509522 371515
rect 509522 371484 509531 371515
rect 509445 371287 509454 371318
rect 509454 371287 509522 371318
rect 509522 371287 509531 371318
rect 509445 371260 509531 371287
rect 509439 370930 509533 370990
rect 52640 359406 53366 360230
rect 142640 359406 143366 360230
rect 232640 359406 233366 360230
rect 322640 359406 323366 360230
rect 417238 368220 417838 368820
rect 420958 368220 421558 368820
rect 412640 359406 413366 360230
rect 507238 368220 507838 368820
rect 510958 368220 511558 368820
rect 502640 359406 503366 360230
rect 64790 263970 65516 264794
rect 57298 254800 57898 255400
rect 61018 254800 61618 255400
rect 153914 263766 154640 264590
rect 146422 254596 147022 255196
rect 150142 254596 150742 255196
rect 245168 263578 245894 264402
rect 334790 263970 335516 264794
rect 424790 263970 425516 264794
rect 514790 263970 515516 264794
rect 58178 251900 58338 252060
rect 234286 252986 234394 253110
rect 149132 252124 149204 252188
rect 59441 251784 59535 251844
rect 60378 251900 60538 252060
rect 59445 251515 59531 251542
rect 59445 251484 59454 251515
rect 59454 251484 59522 251515
rect 59522 251484 59531 251515
rect 59445 251287 59454 251318
rect 59454 251287 59522 251318
rect 59522 251287 59531 251318
rect 59445 251260 59531 251287
rect 147120 251480 147270 251582
rect 149132 251639 149200 251668
rect 149132 251612 149199 251639
rect 149199 251612 149200 251639
rect 149132 251411 149199 251438
rect 149199 251411 149200 251438
rect 149132 251382 149200 251411
rect 232171 251636 232497 251962
rect 151820 251434 151968 251582
rect 234274 251108 234342 251164
rect 59439 250930 59533 250990
rect 149136 251002 149208 251066
rect 57238 248220 57838 248820
rect 249238 250972 249378 251218
rect 320433 251842 321381 252790
rect 329461 250939 329521 250999
rect 329196 250684 329261 250739
rect 60958 248220 61558 248820
rect 52640 239406 53366 240230
rect 146362 248016 146962 248616
rect 150082 248016 150682 248616
rect 141764 239202 142490 240026
rect 337591 248633 339092 250134
rect 420104 251535 420164 251595
rect 419839 251280 419904 251335
rect 411258 248640 412348 249730
rect 233018 239014 233744 239838
rect 428318 249730 429188 250600
rect 510104 251535 510164 251595
rect 509839 251280 509904 251335
rect 501258 248640 502348 249730
rect 518318 249730 519188 250600
rect 322640 239406 323366 240230
rect 412640 239406 413366 240230
rect 502640 239406 503366 240230
rect 57298 148700 57898 149300
rect 61018 148700 61618 149300
rect 147298 148700 147898 149300
rect 151018 148700 151618 149300
rect 237298 148700 237898 149300
rect 241018 148700 241618 149300
rect 327298 148700 327898 149300
rect 331018 148700 331618 149300
rect 417298 148700 417898 149300
rect 421018 148700 421618 149300
rect 507298 148700 507898 149300
rect 511018 148700 511618 149300
rect 58178 145800 58338 145960
rect 60378 145800 60538 145960
rect 148178 145800 148338 145960
rect 150378 145800 150538 145960
rect 238178 145800 238338 145960
rect 240378 145800 240538 145960
rect 328178 145800 328338 145960
rect 330378 145800 330538 145960
rect 418178 145800 418338 145960
rect 420378 145800 420538 145960
rect 508178 145800 508338 145960
rect 510378 145800 510538 145960
rect 57238 142120 57838 142720
rect 60958 142120 61558 142720
rect 147238 142120 147838 142720
rect 150958 142120 151558 142720
rect 237238 142120 237838 142720
rect 240958 142120 241558 142720
rect 327238 142120 327838 142720
rect 330958 142120 331558 142720
rect 417238 142120 417838 142720
rect 420958 142120 421558 142720
rect 507238 142120 507838 142720
rect 510958 142120 511558 142720
rect 57298 58700 57898 59300
rect 61018 58700 61618 59300
rect 147298 58700 147898 59300
rect 151018 58700 151618 59300
rect 237298 58700 237898 59300
rect 241018 58700 241618 59300
rect 327298 58700 327898 59300
rect 331018 58700 331618 59300
rect 417298 58700 417898 59300
rect 421018 58700 421618 59300
rect 507298 58700 507898 59300
rect 511018 58700 511618 59300
rect 58178 55800 58338 55960
rect 60378 55800 60538 55960
rect 148178 55800 148338 55960
rect 150378 55800 150538 55960
rect 238178 55800 238338 55960
rect 240378 55800 240538 55960
rect 328178 55800 328338 55960
rect 330378 55800 330538 55960
rect 418178 55800 418338 55960
rect 420378 55800 420538 55960
rect 508178 55800 508338 55960
rect 510378 55800 510538 55960
rect 57238 52120 57838 52720
rect 60958 52120 61558 52720
rect 147238 52120 147838 52720
rect 150958 52120 151558 52720
rect 237238 52120 237838 52720
rect 240958 52120 241558 52720
rect 327238 52120 327838 52720
rect 330958 52120 331558 52720
rect 417238 52120 417838 52720
rect 420958 52120 421558 52720
rect 507238 52120 507838 52720
rect 510958 52120 511558 52720
<< metal2 >>
rect 326940 664204 327900 664324
rect 326940 663544 327120 664204
rect 327780 663544 327900 664204
rect 57138 662280 58098 662400
rect 57138 661620 57318 662280
rect 57978 661620 58098 662280
rect 57138 659300 58098 661620
rect 57138 658700 57298 659300
rect 57898 658700 58098 659300
rect 60858 662280 61818 662400
rect 60858 661620 61038 662280
rect 61698 661620 61818 662280
rect 60858 659300 61818 661620
rect 60858 658700 61018 659300
rect 61618 658700 61818 659300
rect 147138 662280 148098 662400
rect 147138 661620 147318 662280
rect 147978 661620 148098 662280
rect 147138 659300 148098 661620
rect 147138 658700 147298 659300
rect 147898 658700 148098 659300
rect 150858 662280 151818 662400
rect 150858 661620 151038 662280
rect 151698 661620 151818 662280
rect 150858 659300 151818 661620
rect 150858 658700 151018 659300
rect 151618 658700 151818 659300
rect 237138 662280 238098 662400
rect 237138 661620 237318 662280
rect 237978 661620 238098 662280
rect 237138 659300 238098 661620
rect 237138 658700 237298 659300
rect 237898 658700 238098 659300
rect 240858 662280 241818 662400
rect 240858 661620 241038 662280
rect 241698 661620 241818 662280
rect 240858 659300 241818 661620
rect 326940 661224 327900 663544
rect 326940 660624 327100 661224
rect 327700 660624 327900 661224
rect 330660 664204 331620 664324
rect 330660 663544 330840 664204
rect 331500 663544 331620 664204
rect 330660 661224 331620 663544
rect 330660 660624 330820 661224
rect 331420 660624 331620 661224
rect 416940 664204 417900 664324
rect 416940 663544 417120 664204
rect 417780 663544 417900 664204
rect 416940 661224 417900 663544
rect 416940 660624 417100 661224
rect 417700 660624 417900 661224
rect 420660 664204 421620 664324
rect 420660 663544 420840 664204
rect 421500 663544 421620 664204
rect 420660 661224 421620 663544
rect 420660 660624 420820 661224
rect 421420 660624 421620 661224
rect 506940 664204 507900 664324
rect 506940 663544 507120 664204
rect 507780 663544 507900 664204
rect 506940 661224 507900 663544
rect 506940 660624 507100 661224
rect 507700 660624 507900 661224
rect 510660 664204 511620 664324
rect 510660 663544 510840 664204
rect 511500 663544 511620 664204
rect 510660 661224 511620 663544
rect 510660 660624 510820 661224
rect 511420 660624 511620 661224
rect 240858 658700 241018 659300
rect 241618 658700 241818 659300
rect 327960 657884 328160 657904
rect 327960 657724 327980 657884
rect 328140 657724 328160 657884
rect 327960 657124 328160 657724
rect 330160 657884 330360 657904
rect 330160 657724 330180 657884
rect 330340 657864 330360 657884
rect 417960 657884 418160 657904
rect 330340 657854 330440 657864
rect 330340 657754 330890 657854
rect 330340 657744 330440 657754
rect 330340 657724 330360 657744
rect 330160 657704 330360 657724
rect 330790 657734 330890 657754
rect 331440 657764 331640 657784
rect 331440 657734 331460 657764
rect 330790 657634 331460 657734
rect 331440 657604 331460 657634
rect 331620 657604 331640 657764
rect 331440 657584 331640 657604
rect 417960 657724 417980 657884
rect 418140 657724 418160 657884
rect 417960 657124 418160 657724
rect 420160 657884 420360 657904
rect 420160 657724 420180 657884
rect 420340 657864 420360 657884
rect 507960 657884 508160 657904
rect 420340 657854 420440 657864
rect 420340 657754 420890 657854
rect 420340 657744 420440 657754
rect 420340 657724 420360 657744
rect 420160 657704 420360 657724
rect 420790 657734 420890 657754
rect 421440 657764 421640 657784
rect 421440 657734 421460 657764
rect 420790 657634 421460 657734
rect 421440 657604 421460 657634
rect 421620 657604 421640 657764
rect 421440 657584 421640 657604
rect 507960 657724 507980 657884
rect 508140 657724 508160 657884
rect 507960 657124 508160 657724
rect 510160 657884 510360 657904
rect 510160 657724 510180 657884
rect 510340 657864 510360 657884
rect 510340 657854 510440 657864
rect 510340 657754 510890 657854
rect 510340 657744 510440 657754
rect 510340 657724 510360 657744
rect 510160 657704 510360 657724
rect 510790 657734 510890 657754
rect 511440 657764 511640 657784
rect 511440 657734 511460 657764
rect 510790 657634 511460 657734
rect 511440 657604 511460 657634
rect 511620 657604 511640 657764
rect 511440 657584 511640 657604
rect 327320 657084 328160 657124
rect 327320 656964 327360 657084
rect 327560 656964 328160 657084
rect 327320 656924 328160 656964
rect 417320 657084 418160 657124
rect 417320 656964 417360 657084
rect 417560 656964 418160 657084
rect 417320 656924 418160 656964
rect 507320 657084 508160 657124
rect 507320 656964 507360 657084
rect 507560 656964 508160 657084
rect 507320 656924 508160 656964
rect 58158 655960 58358 655980
rect 58158 655800 58178 655960
rect 58338 655800 58358 655960
rect 58158 655200 58358 655800
rect 60358 655960 60558 655980
rect 60358 655800 60378 655960
rect 60538 655940 60558 655960
rect 148158 655960 148358 655980
rect 60538 655930 60638 655940
rect 60538 655830 61088 655930
rect 60538 655820 60638 655830
rect 60538 655800 60558 655820
rect 60358 655780 60558 655800
rect 60988 655810 61088 655830
rect 61638 655840 61838 655860
rect 61638 655810 61658 655840
rect 60988 655710 61658 655810
rect 61638 655680 61658 655710
rect 61818 655680 61838 655840
rect 61638 655660 61838 655680
rect 148158 655800 148178 655960
rect 148338 655800 148358 655960
rect 148158 655200 148358 655800
rect 150358 655960 150558 655980
rect 150358 655800 150378 655960
rect 150538 655940 150558 655960
rect 238158 655960 238358 655980
rect 150538 655930 150638 655940
rect 150538 655830 151088 655930
rect 150538 655820 150638 655830
rect 150538 655800 150558 655820
rect 150358 655780 150558 655800
rect 150988 655810 151088 655830
rect 151638 655840 151838 655860
rect 151638 655810 151658 655840
rect 150988 655710 151658 655810
rect 151638 655680 151658 655710
rect 151818 655680 151838 655840
rect 151638 655660 151838 655680
rect 238158 655800 238178 655960
rect 238338 655800 238358 655960
rect 238158 655200 238358 655800
rect 240358 655960 240558 655980
rect 240358 655800 240378 655960
rect 240538 655940 240558 655960
rect 240538 655930 240638 655940
rect 240538 655830 241088 655930
rect 240538 655820 240638 655830
rect 240538 655800 240558 655820
rect 240358 655780 240558 655800
rect 240988 655810 241088 655830
rect 241638 655840 241838 655860
rect 241638 655810 241658 655840
rect 240988 655710 241658 655810
rect 241638 655680 241658 655710
rect 241818 655680 241838 655840
rect 241638 655660 241838 655680
rect 57518 655160 58358 655200
rect 57518 655040 57558 655160
rect 57758 655040 58358 655160
rect 57518 655000 58358 655040
rect 147518 655160 148358 655200
rect 147518 655040 147558 655160
rect 147758 655040 148358 655160
rect 147518 655000 148358 655040
rect 237518 655160 238358 655200
rect 237518 655040 237558 655160
rect 237758 655040 238358 655160
rect 237518 655000 238358 655040
rect 326880 654044 327040 654644
rect 327640 654044 327840 654644
rect 57078 652120 57238 652720
rect 57838 652120 58038 652720
rect 57078 649800 58038 652120
rect 57078 649140 57258 649800
rect 57918 649140 58038 649800
rect 57078 649020 58038 649140
rect 60798 652120 60958 652720
rect 61558 652120 61758 652720
rect 60798 649800 61758 652120
rect 60798 649140 60978 649800
rect 61638 649140 61758 649800
rect 60798 649020 61758 649140
rect 147078 652120 147238 652720
rect 147838 652120 148038 652720
rect 147078 649800 148038 652120
rect 147078 649140 147258 649800
rect 147918 649140 148038 649800
rect 147078 649020 148038 649140
rect 150798 652120 150958 652720
rect 151558 652120 151758 652720
rect 150798 649800 151758 652120
rect 150798 649140 150978 649800
rect 151638 649140 151758 649800
rect 150798 649020 151758 649140
rect 237078 652120 237238 652720
rect 237838 652120 238038 652720
rect 237078 649800 238038 652120
rect 237078 649140 237258 649800
rect 237918 649140 238038 649800
rect 237078 649020 238038 649140
rect 240798 652120 240958 652720
rect 241558 652120 241758 652720
rect 240798 649800 241758 652120
rect 326880 651724 327840 654044
rect 326880 651064 327060 651724
rect 327720 651064 327840 651724
rect 326880 650944 327840 651064
rect 330600 654044 330760 654644
rect 331360 654044 331560 654644
rect 330600 651724 331560 654044
rect 330600 651064 330780 651724
rect 331440 651064 331560 651724
rect 330600 650944 331560 651064
rect 416880 654044 417040 654644
rect 417640 654044 417840 654644
rect 416880 651724 417840 654044
rect 416880 651064 417060 651724
rect 417720 651064 417840 651724
rect 416880 650944 417840 651064
rect 420600 654044 420760 654644
rect 421360 654044 421560 654644
rect 420600 651724 421560 654044
rect 420600 651064 420780 651724
rect 421440 651064 421560 651724
rect 420600 650944 421560 651064
rect 506880 654044 507040 654644
rect 507640 654044 507840 654644
rect 506880 651724 507840 654044
rect 506880 651064 507060 651724
rect 507720 651064 507840 651724
rect 506880 650944 507840 651064
rect 510600 654044 510760 654644
rect 511360 654044 511560 654644
rect 510600 651724 511560 654044
rect 510600 651064 510780 651724
rect 511440 651064 511560 651724
rect 510600 650944 511560 651064
rect 240798 649140 240978 649800
rect 241638 649140 241758 649800
rect 240798 649020 241758 649140
rect 416940 589204 417900 589324
rect 416940 588544 417120 589204
rect 417780 588544 417900 589204
rect 57138 587280 58098 587400
rect 57138 586620 57318 587280
rect 57978 586620 58098 587280
rect 57138 584300 58098 586620
rect 57138 583700 57298 584300
rect 57898 583700 58098 584300
rect 60858 587280 61818 587400
rect 60858 586620 61038 587280
rect 61698 586620 61818 587280
rect 60858 584300 61818 586620
rect 60858 583700 61018 584300
rect 61618 583700 61818 584300
rect 147138 587280 148098 587400
rect 147138 586620 147318 587280
rect 147978 586620 148098 587280
rect 147138 584300 148098 586620
rect 147138 583700 147298 584300
rect 147898 583700 148098 584300
rect 150858 587280 151818 587400
rect 150858 586620 151038 587280
rect 151698 586620 151818 587280
rect 150858 584300 151818 586620
rect 150858 583700 151018 584300
rect 151618 583700 151818 584300
rect 237138 587280 238098 587400
rect 237138 586620 237318 587280
rect 237978 586620 238098 587280
rect 237138 584300 238098 586620
rect 237138 583700 237298 584300
rect 237898 583700 238098 584300
rect 240858 587280 241818 587400
rect 240858 586620 241038 587280
rect 241698 586620 241818 587280
rect 240858 584300 241818 586620
rect 240858 583700 241018 584300
rect 241618 583700 241818 584300
rect 327138 587280 328098 587400
rect 327138 586620 327318 587280
rect 327978 586620 328098 587280
rect 327138 584300 328098 586620
rect 327138 583700 327298 584300
rect 327898 583700 328098 584300
rect 330858 587280 331818 587400
rect 330858 586620 331038 587280
rect 331698 586620 331818 587280
rect 330858 584300 331818 586620
rect 416940 586224 417900 588544
rect 416940 585624 417100 586224
rect 417700 585624 417900 586224
rect 420660 589204 421620 589324
rect 420660 588544 420840 589204
rect 421500 588544 421620 589204
rect 420660 586224 421620 588544
rect 420660 585624 420820 586224
rect 421420 585624 421620 586224
rect 506940 589204 507900 589324
rect 506940 588544 507120 589204
rect 507780 588544 507900 589204
rect 506940 586224 507900 588544
rect 506940 585624 507100 586224
rect 507700 585624 507900 586224
rect 510660 589204 511620 589324
rect 510660 588544 510840 589204
rect 511500 588544 511620 589204
rect 510660 586224 511620 588544
rect 510660 585624 510820 586224
rect 511420 585624 511620 586224
rect 330858 583700 331018 584300
rect 331618 583700 331818 584300
rect 417960 582884 418160 582904
rect 417960 582724 417980 582884
rect 418140 582724 418160 582884
rect 417960 582124 418160 582724
rect 420160 582884 420360 582904
rect 420160 582724 420180 582884
rect 420340 582864 420360 582884
rect 507960 582884 508160 582904
rect 420340 582854 420440 582864
rect 420340 582754 420890 582854
rect 420340 582744 420440 582754
rect 420340 582724 420360 582744
rect 420160 582704 420360 582724
rect 420790 582734 420890 582754
rect 421440 582764 421640 582784
rect 421440 582734 421460 582764
rect 420790 582634 421460 582734
rect 421440 582604 421460 582634
rect 421620 582604 421640 582764
rect 421440 582584 421640 582604
rect 507960 582724 507980 582884
rect 508140 582724 508160 582884
rect 507960 582124 508160 582724
rect 510160 582884 510360 582904
rect 510160 582724 510180 582884
rect 510340 582864 510360 582884
rect 510340 582854 510440 582864
rect 510340 582754 510890 582854
rect 510340 582744 510440 582754
rect 510340 582724 510360 582744
rect 510160 582704 510360 582724
rect 510790 582734 510890 582754
rect 511440 582764 511640 582784
rect 511440 582734 511460 582764
rect 510790 582634 511460 582734
rect 511440 582604 511460 582634
rect 511620 582604 511640 582764
rect 511440 582584 511640 582604
rect 417320 582084 418160 582124
rect 417320 581964 417360 582084
rect 417560 581964 418160 582084
rect 417320 581924 418160 581964
rect 507320 582084 508160 582124
rect 507320 581964 507360 582084
rect 507560 581964 508160 582084
rect 507320 581924 508160 581964
rect 58158 580960 58358 580980
rect 58158 580800 58178 580960
rect 58338 580800 58358 580960
rect 58158 580200 58358 580800
rect 60358 580960 60558 580980
rect 60358 580800 60378 580960
rect 60538 580940 60558 580960
rect 148158 580960 148358 580980
rect 60538 580930 60638 580940
rect 60538 580830 61088 580930
rect 60538 580820 60638 580830
rect 60538 580800 60558 580820
rect 60358 580780 60558 580800
rect 60988 580810 61088 580830
rect 61638 580840 61838 580860
rect 61638 580810 61658 580840
rect 60988 580710 61658 580810
rect 61638 580680 61658 580710
rect 61818 580680 61838 580840
rect 61638 580660 61838 580680
rect 148158 580800 148178 580960
rect 148338 580800 148358 580960
rect 148158 580200 148358 580800
rect 150358 580960 150558 580980
rect 150358 580800 150378 580960
rect 150538 580940 150558 580960
rect 238158 580960 238358 580980
rect 150538 580930 150638 580940
rect 150538 580830 151088 580930
rect 150538 580820 150638 580830
rect 150538 580800 150558 580820
rect 150358 580780 150558 580800
rect 150988 580810 151088 580830
rect 151638 580840 151838 580860
rect 151638 580810 151658 580840
rect 150988 580710 151658 580810
rect 151638 580680 151658 580710
rect 151818 580680 151838 580840
rect 151638 580660 151838 580680
rect 238158 580800 238178 580960
rect 238338 580800 238358 580960
rect 238158 580200 238358 580800
rect 240358 580960 240558 580980
rect 240358 580800 240378 580960
rect 240538 580940 240558 580960
rect 328158 580960 328358 580980
rect 240538 580930 240638 580940
rect 240538 580830 241088 580930
rect 240538 580820 240638 580830
rect 240538 580800 240558 580820
rect 240358 580780 240558 580800
rect 240988 580810 241088 580830
rect 241638 580840 241838 580860
rect 241638 580810 241658 580840
rect 240988 580710 241658 580810
rect 241638 580680 241658 580710
rect 241818 580680 241838 580840
rect 241638 580660 241838 580680
rect 328158 580800 328178 580960
rect 328338 580800 328358 580960
rect 328158 580200 328358 580800
rect 330358 580960 330558 580980
rect 330358 580800 330378 580960
rect 330538 580940 330558 580960
rect 330538 580930 330638 580940
rect 330538 580830 331088 580930
rect 330538 580820 330638 580830
rect 330538 580800 330558 580820
rect 330358 580780 330558 580800
rect 330988 580810 331088 580830
rect 331638 580840 331838 580860
rect 331638 580810 331658 580840
rect 330988 580710 331658 580810
rect 331638 580680 331658 580710
rect 331818 580680 331838 580840
rect 331638 580660 331838 580680
rect 57518 580160 58358 580200
rect 57518 580040 57558 580160
rect 57758 580040 58358 580160
rect 57518 580000 58358 580040
rect 147518 580160 148358 580200
rect 147518 580040 147558 580160
rect 147758 580040 148358 580160
rect 147518 580000 148358 580040
rect 237518 580160 238358 580200
rect 237518 580040 237558 580160
rect 237758 580040 238358 580160
rect 237518 580000 238358 580040
rect 327518 580160 328358 580200
rect 327518 580040 327558 580160
rect 327758 580040 328358 580160
rect 327518 580000 328358 580040
rect 416880 579044 417040 579644
rect 417640 579044 417840 579644
rect 57078 577120 57238 577720
rect 57838 577120 58038 577720
rect 57078 574800 58038 577120
rect 57078 574140 57258 574800
rect 57918 574140 58038 574800
rect 57078 574020 58038 574140
rect 60798 577120 60958 577720
rect 61558 577120 61758 577720
rect 60798 574800 61758 577120
rect 60798 574140 60978 574800
rect 61638 574140 61758 574800
rect 60798 574020 61758 574140
rect 147078 577120 147238 577720
rect 147838 577120 148038 577720
rect 147078 574800 148038 577120
rect 147078 574140 147258 574800
rect 147918 574140 148038 574800
rect 147078 574020 148038 574140
rect 150798 577120 150958 577720
rect 151558 577120 151758 577720
rect 150798 574800 151758 577120
rect 150798 574140 150978 574800
rect 151638 574140 151758 574800
rect 150798 574020 151758 574140
rect 237078 577120 237238 577720
rect 237838 577120 238038 577720
rect 237078 574800 238038 577120
rect 237078 574140 237258 574800
rect 237918 574140 238038 574800
rect 237078 574020 238038 574140
rect 240798 577120 240958 577720
rect 241558 577120 241758 577720
rect 240798 574800 241758 577120
rect 240798 574140 240978 574800
rect 241638 574140 241758 574800
rect 240798 574020 241758 574140
rect 327078 577120 327238 577720
rect 327838 577120 328038 577720
rect 327078 574800 328038 577120
rect 327078 574140 327258 574800
rect 327918 574140 328038 574800
rect 327078 574020 328038 574140
rect 330798 577120 330958 577720
rect 331558 577120 331758 577720
rect 330798 574800 331758 577120
rect 416880 576724 417840 579044
rect 416880 576064 417060 576724
rect 417720 576064 417840 576724
rect 416880 575944 417840 576064
rect 420600 579044 420760 579644
rect 421360 579044 421560 579644
rect 420600 576724 421560 579044
rect 420600 576064 420780 576724
rect 421440 576064 421560 576724
rect 420600 575944 421560 576064
rect 506880 579044 507040 579644
rect 507640 579044 507840 579644
rect 506880 576724 507840 579044
rect 506880 576064 507060 576724
rect 507720 576064 507840 576724
rect 506880 575944 507840 576064
rect 510600 579044 510760 579644
rect 511360 579044 511560 579644
rect 510600 576724 511560 579044
rect 510600 576064 510780 576724
rect 511440 576064 511560 576724
rect 510600 575944 511560 576064
rect 330798 574140 330978 574800
rect 331638 574140 331758 574800
rect 330798 574020 331758 574140
rect 64428 506810 65748 507240
rect 64428 506084 64790 506810
rect 65482 506084 65748 506810
rect 64428 504794 65748 506084
rect 64428 503970 64790 504794
rect 65516 503970 65748 504794
rect 64428 503608 65748 503970
rect 154428 506810 155748 507240
rect 154428 506084 154790 506810
rect 155482 506084 155748 506810
rect 154428 504794 155748 506084
rect 154428 503970 154790 504794
rect 155516 503970 155748 504794
rect 154428 503608 155748 503970
rect 244428 506810 245748 507240
rect 244428 506084 244790 506810
rect 245482 506084 245748 506810
rect 244428 504794 245748 506084
rect 244428 503970 244790 504794
rect 245516 503970 245748 504794
rect 244428 503608 245748 503970
rect 334428 506810 335748 507240
rect 334428 506084 334790 506810
rect 335482 506084 335748 506810
rect 334428 504794 335748 506084
rect 334428 503970 334790 504794
rect 335516 503970 335748 504794
rect 334428 503608 335748 503970
rect 424428 506810 425748 507240
rect 424428 506084 424790 506810
rect 425482 506084 425748 506810
rect 424428 504794 425748 506084
rect 424428 503970 424790 504794
rect 425516 503970 425748 504794
rect 424428 503608 425748 503970
rect 514428 506810 515748 507240
rect 514428 506084 514790 506810
rect 515482 506084 515748 506810
rect 514428 504794 515748 506084
rect 514428 503970 514790 504794
rect 515516 503970 515748 504794
rect 514428 503608 515748 503970
rect 147108 499935 148093 500105
rect 147108 499190 147278 499935
rect 147958 499190 148093 499935
rect 147108 498510 148093 499190
rect 150828 499965 151828 500055
rect 150828 499220 150998 499965
rect 151678 499220 151828 499965
rect 57138 498380 58098 498500
rect 57138 497720 57318 498380
rect 57978 497720 58098 498380
rect 57138 495400 58098 497720
rect 57138 494800 57298 495400
rect 57898 494800 58098 495400
rect 60858 498380 61818 498500
rect 60858 497720 61038 498380
rect 61698 497720 61818 498380
rect 60858 495400 61818 497720
rect 147433 496895 147633 498510
rect 150828 498460 151828 499220
rect 151203 496895 151403 498460
rect 147433 496695 151403 496895
rect 237138 498380 238098 498500
rect 237138 497720 237318 498380
rect 237978 497720 238098 498380
rect 60858 494800 61018 495400
rect 61618 494800 61818 495400
rect 60000 492392 60086 492401
rect 60000 492328 60008 492392
rect 60080 492328 60086 492392
rect 60000 491872 60086 492328
rect 150039 492200 150239 496695
rect 237138 495843 238098 497720
rect 240858 498380 241818 498500
rect 240858 497720 241038 498380
rect 241698 497720 241818 498380
rect 240858 495843 241818 497720
rect 327138 498380 328098 498500
rect 327138 497720 327318 498380
rect 327978 497720 328098 498380
rect 327138 496829 328098 497720
rect 330858 498380 331818 498500
rect 330858 497720 331038 498380
rect 331698 497720 331818 498380
rect 330858 496829 331818 497720
rect 417138 498380 418098 498500
rect 417138 497720 417318 498380
rect 417978 497720 418098 498380
rect 324728 496814 331827 496829
rect 237086 495282 241819 495843
rect 323734 495757 331827 496814
rect 237138 495278 238098 495282
rect 230424 493495 230433 494443
rect 231381 493495 231390 494443
rect 230433 492790 231381 493495
rect 57544 491794 58162 491830
rect 60000 491816 60008 491872
rect 60076 491816 60086 491872
rect 60000 491808 60086 491816
rect 57544 491668 57598 491794
rect 57746 491786 58162 491794
rect 57746 491684 57996 491786
rect 58146 491684 58162 491786
rect 57746 491668 58162 491684
rect 57544 491638 58162 491668
rect 62664 491786 62866 491814
rect 60000 491642 60086 491650
rect 60000 491586 60008 491642
rect 60076 491586 60086 491642
rect 60000 491270 60086 491586
rect 60000 491206 60012 491270
rect 60084 491206 60086 491270
rect 60000 491189 60086 491206
rect 62664 491638 62696 491786
rect 62844 491638 62866 491786
rect 62664 491408 62866 491638
rect 150094 491595 150189 492200
rect 230427 491842 230433 492790
rect 231381 491842 231387 492790
rect 239396 491604 239596 495282
rect 240858 495261 241818 495282
rect 323734 493596 324296 495757
rect 417138 495400 418098 497720
rect 417138 494800 417298 495400
rect 417898 494800 418098 495400
rect 420858 498380 421818 498500
rect 420858 497720 421038 498380
rect 421698 497720 421818 498380
rect 420858 495400 421818 497720
rect 420858 494800 421018 495400
rect 421618 494800 421818 495400
rect 507138 498380 508098 498500
rect 507138 497720 507318 498380
rect 507978 497720 508098 498380
rect 507138 495400 508098 497720
rect 507138 494800 507298 495400
rect 507898 494800 508098 495400
rect 510858 498380 511818 498500
rect 510858 497720 511038 498380
rect 511698 497720 511818 498380
rect 510858 495400 511818 497720
rect 510858 494800 511018 495400
rect 511618 494800 511818 495400
rect 323744 493502 324280 493596
rect 323744 493378 323908 493502
rect 324016 493378 324280 493502
rect 323744 493216 324280 493378
rect 510000 492392 510086 492401
rect 321793 492354 322119 492360
rect 320954 492028 320963 492354
rect 321289 492028 321793 492354
rect 510000 492328 510008 492392
rect 510080 492328 510086 492392
rect 321793 492022 322119 492028
rect 418158 492060 418358 492080
rect 418158 491900 418178 492060
rect 418338 491900 418358 492060
rect 338796 491700 339592 491702
rect 338796 491610 339791 491700
rect 150094 491535 150104 491595
rect 150164 491535 150189 491595
rect 150094 491525 150189 491535
rect 62664 491204 62700 491408
rect 62830 491204 62866 491408
rect 62664 491178 62866 491204
rect 149829 491335 149914 491340
rect 149829 491280 149839 491335
rect 149904 491280 149914 491335
rect 149829 491265 149914 491280
rect 149829 490350 149911 491265
rect 239451 490999 239546 491604
rect 239451 490939 239461 490999
rect 239521 490939 239546 490999
rect 239451 490929 239546 490939
rect 323888 491556 323970 491574
rect 323888 491500 323896 491556
rect 323964 491500 323970 491556
rect 239186 490739 239271 490744
rect 239186 490684 239196 490739
rect 239261 490684 239271 490739
rect 239186 490669 239271 490684
rect 57078 488220 57238 488820
rect 57838 488220 58038 488820
rect 57078 485900 58038 488220
rect 57078 485240 57258 485900
rect 57918 485240 58038 485900
rect 57078 485120 58038 485240
rect 60798 488220 60958 488820
rect 61558 488220 61758 488820
rect 139654 488640 139663 489730
rect 140753 488640 141258 489730
rect 142348 488640 142354 489730
rect 149769 489630 149979 490350
rect 158312 489730 158318 490600
rect 159188 489730 159194 490600
rect 239186 489754 239268 490669
rect 323888 490326 323970 491500
rect 338796 491364 338860 491610
rect 339000 491364 339791 491610
rect 338796 491282 339791 491364
rect 339192 491278 339791 491282
rect 340213 491278 340222 491700
rect 418158 491300 418358 491900
rect 420358 492060 420558 492080
rect 420358 491900 420378 492060
rect 420538 492040 420558 492060
rect 420538 492030 420638 492040
rect 420538 491930 421088 492030
rect 420538 491920 420638 491930
rect 420538 491900 420558 491920
rect 420358 491880 420558 491900
rect 420988 491910 421088 491930
rect 421638 491940 421838 491960
rect 421638 491910 421658 491940
rect 419401 491844 419573 491864
rect 419401 491784 419441 491844
rect 419535 491784 419573 491844
rect 420988 491810 421658 491910
rect 419401 491756 419573 491784
rect 421638 491780 421658 491810
rect 421818 491780 421838 491940
rect 510000 491872 510086 492328
rect 421638 491760 421838 491780
rect 507544 491794 508162 491830
rect 510000 491816 510008 491872
rect 510076 491816 510086 491872
rect 510000 491808 510086 491816
rect 419437 491542 419539 491756
rect 507544 491668 507598 491794
rect 507746 491786 508162 491794
rect 507746 491684 507996 491786
rect 508146 491684 508162 491786
rect 507746 491668 508162 491684
rect 507544 491638 508162 491668
rect 512664 491786 512866 491814
rect 510000 491642 510086 491650
rect 419437 491484 419445 491542
rect 419531 491484 419539 491542
rect 419437 491478 419539 491484
rect 510000 491586 510008 491642
rect 510076 491586 510086 491642
rect 417518 491260 418358 491300
rect 417518 491140 417558 491260
rect 417758 491140 418358 491260
rect 417518 491100 418358 491140
rect 419437 491318 419539 491322
rect 419437 491260 419445 491318
rect 419531 491260 419539 491318
rect 419437 491014 419539 491260
rect 510000 491270 510086 491586
rect 510000 491206 510012 491270
rect 510084 491206 510086 491270
rect 510000 491189 510086 491206
rect 512664 491638 512696 491786
rect 512844 491638 512866 491786
rect 512664 491408 512866 491638
rect 512664 491204 512700 491408
rect 512830 491204 512866 491408
rect 512664 491178 512866 491204
rect 419397 490990 419569 491014
rect 419397 490930 419439 490990
rect 419533 490930 419569 490990
rect 419397 490906 419569 490930
rect 330798 490326 331758 490328
rect 147478 489420 151438 489630
rect 60798 485900 61758 488220
rect 147478 486940 147688 489420
rect 151228 486965 151438 489420
rect 158318 489300 159188 489730
rect 158318 488421 159188 488430
rect 237088 488517 238038 488525
rect 239126 488517 239336 489754
rect 247585 488633 247591 490134
rect 249092 488633 249098 490134
rect 323880 489374 331774 490326
rect 240798 488517 241743 488547
rect 237088 488178 241743 488517
rect 237088 488000 238038 488178
rect 60798 485240 60978 485900
rect 61638 485240 61758 485900
rect 60798 485120 61758 485240
rect 147038 485130 148073 486940
rect 147038 484385 147193 485130
rect 147873 484385 148073 485130
rect 150793 485130 151758 486965
rect 150793 484385 150963 485130
rect 151643 484385 151758 485130
rect 237078 485900 238038 488000
rect 237078 485240 237258 485900
rect 237918 485240 238038 485900
rect 237078 485120 238038 485240
rect 240798 487812 241743 488178
rect 247591 488088 249092 488633
rect 240798 485900 241758 487812
rect 247591 486578 249092 486587
rect 240798 485240 240978 485900
rect 241638 485240 241758 485900
rect 240798 485120 241758 485240
rect 327078 485900 328038 489374
rect 327078 485240 327258 485900
rect 327918 485240 328038 485900
rect 327078 485120 328038 485240
rect 330798 485900 331758 489374
rect 330798 485240 330978 485900
rect 331638 485240 331758 485900
rect 330798 485120 331758 485240
rect 417078 488220 417238 488820
rect 417838 488220 418038 488820
rect 417078 485900 418038 488220
rect 417078 485240 417258 485900
rect 417918 485240 418038 485900
rect 417078 485120 418038 485240
rect 420798 488220 420958 488820
rect 421558 488220 421758 488820
rect 420798 485900 421758 488220
rect 420798 485240 420978 485900
rect 421638 485240 421758 485900
rect 420798 485120 421758 485240
rect 507078 488220 507238 488820
rect 507838 488220 508038 488820
rect 507078 485900 508038 488220
rect 507078 485240 507258 485900
rect 507918 485240 508038 485900
rect 507078 485120 508038 485240
rect 510798 488220 510958 488820
rect 511558 488220 511758 488820
rect 510798 485900 511758 488220
rect 510798 485240 510978 485900
rect 511638 485240 511758 485900
rect 510798 485120 511758 485240
rect 147038 484275 148073 484385
rect 52344 480230 53664 480398
rect 52344 479406 52640 480230
rect 53366 479406 53664 480230
rect 52344 477788 53664 479406
rect 52344 477062 52608 477788
rect 53300 477062 53664 477788
rect 52344 476766 53664 477062
rect 142344 480230 143664 480398
rect 142344 479406 142640 480230
rect 143366 479406 143664 480230
rect 142344 477788 143664 479406
rect 142344 477062 142608 477788
rect 143300 477062 143664 477788
rect 142344 476766 143664 477062
rect 232344 480230 233664 480398
rect 232344 479406 232640 480230
rect 233366 479406 233664 480230
rect 232344 477788 233664 479406
rect 232344 477062 232608 477788
rect 233300 477062 233664 477788
rect 232344 476766 233664 477062
rect 322344 480230 323664 480398
rect 322344 479406 322640 480230
rect 323366 479406 323664 480230
rect 322344 477788 323664 479406
rect 322344 477062 322608 477788
rect 323300 477062 323664 477788
rect 322344 476766 323664 477062
rect 412344 480230 413664 480398
rect 412344 479406 412640 480230
rect 413366 479406 413664 480230
rect 412344 477788 413664 479406
rect 412344 477062 412608 477788
rect 413300 477062 413664 477788
rect 412344 476766 413664 477062
rect 502344 480230 503664 480398
rect 502344 479406 502640 480230
rect 503366 479406 503664 480230
rect 502344 477788 503664 479406
rect 502344 477062 502608 477788
rect 503300 477062 503664 477788
rect 502344 476766 503664 477062
rect 64428 386810 65748 387240
rect 64428 386084 64790 386810
rect 65482 386084 65748 386810
rect 64428 384794 65748 386084
rect 64428 383970 64790 384794
rect 65516 383970 65748 384794
rect 64428 383608 65748 383970
rect 154428 386810 155748 387240
rect 154428 386084 154790 386810
rect 155482 386084 155748 386810
rect 154428 384794 155748 386084
rect 154428 383970 154790 384794
rect 155516 383970 155748 384794
rect 154428 383608 155748 383970
rect 244428 386810 245748 387240
rect 244428 386084 244790 386810
rect 245482 386084 245748 386810
rect 244428 384794 245748 386084
rect 244428 383970 244790 384794
rect 245516 383970 245748 384794
rect 244428 383608 245748 383970
rect 334428 386810 335748 387240
rect 334428 386084 334790 386810
rect 335482 386084 335748 386810
rect 334428 384794 335748 386084
rect 334428 383970 334790 384794
rect 335516 383970 335748 384794
rect 334428 383608 335748 383970
rect 424428 386810 425748 387240
rect 424428 386084 424790 386810
rect 425482 386084 425748 386810
rect 424428 384794 425748 386084
rect 424428 383970 424790 384794
rect 425516 383970 425748 384794
rect 424428 383608 425748 383970
rect 514428 386810 515748 387240
rect 514428 386084 514790 386810
rect 515482 386084 515748 386810
rect 514428 384794 515748 386084
rect 514428 383970 514790 384794
rect 515516 383970 515748 384794
rect 514428 383608 515748 383970
rect 57108 379935 58093 380105
rect 57108 379190 57278 379935
rect 57958 379190 58093 379935
rect 57108 378510 58093 379190
rect 60828 379965 61828 380055
rect 60828 379220 60998 379965
rect 61678 379220 61828 379965
rect 57433 376895 57633 378510
rect 60828 378460 61828 379220
rect 147108 379935 148093 380105
rect 147108 379190 147278 379935
rect 147958 379190 148093 379935
rect 147108 378510 148093 379190
rect 150828 379965 151828 380055
rect 150828 379220 150998 379965
rect 151678 379220 151828 379965
rect 61203 376895 61403 378460
rect 57433 376695 61403 376895
rect 147433 376895 147633 378510
rect 150828 378460 151828 379220
rect 151203 376895 151403 378460
rect 147433 376695 151403 376895
rect 237138 378380 238098 378500
rect 237138 377720 237318 378380
rect 237978 377720 238098 378380
rect 60039 372200 60239 376695
rect 150039 372200 150239 376695
rect 237138 375843 238098 377720
rect 240858 378380 241818 378500
rect 240858 377720 241038 378380
rect 241698 377720 241818 378380
rect 240858 375843 241818 377720
rect 327138 378380 328098 378500
rect 327138 377720 327318 378380
rect 327978 377720 328098 378380
rect 327138 376829 328098 377720
rect 330858 378380 331818 378500
rect 330858 377720 331038 378380
rect 331698 377720 331818 378380
rect 330858 376829 331818 377720
rect 417138 378380 418098 378500
rect 417138 377720 417318 378380
rect 417978 377720 418098 378380
rect 324728 376814 331827 376829
rect 237086 375282 241819 375843
rect 323734 375757 331827 376814
rect 237138 375278 238098 375282
rect 230424 373495 230433 374443
rect 231381 373495 231390 374443
rect 230433 372790 231381 373495
rect 60094 371595 60189 372200
rect 60094 371535 60104 371595
rect 60164 371535 60189 371595
rect 60094 371525 60189 371535
rect 150094 371595 150189 372200
rect 230427 371842 230433 372790
rect 231381 371842 231387 372790
rect 239396 371604 239596 375282
rect 240858 375261 241818 375282
rect 323734 373596 324296 375757
rect 417138 375400 418098 377720
rect 417138 374800 417298 375400
rect 417898 374800 418098 375400
rect 420858 378380 421818 378500
rect 420858 377720 421038 378380
rect 421698 377720 421818 378380
rect 420858 375400 421818 377720
rect 420858 374800 421018 375400
rect 421618 374800 421818 375400
rect 507138 378380 508098 378500
rect 507138 377720 507318 378380
rect 507978 377720 508098 378380
rect 507138 375400 508098 377720
rect 507138 374800 507298 375400
rect 507898 374800 508098 375400
rect 510858 378380 511818 378500
rect 510858 377720 511038 378380
rect 511698 377720 511818 378380
rect 510858 375400 511818 377720
rect 510858 374800 511018 375400
rect 511618 374800 511818 375400
rect 323744 373502 324280 373596
rect 323744 373378 323908 373502
rect 324016 373378 324280 373502
rect 323744 373216 324280 373378
rect 420000 372392 420086 372401
rect 321793 372354 322119 372360
rect 320954 372028 320963 372354
rect 321289 372028 321793 372354
rect 321793 372022 322119 372028
rect 420000 372328 420008 372392
rect 420080 372328 420086 372392
rect 420000 371872 420086 372328
rect 417544 371794 418162 371830
rect 420000 371816 420008 371872
rect 420076 371816 420086 371872
rect 420000 371808 420086 371816
rect 508158 372060 508358 372080
rect 508158 371900 508178 372060
rect 508338 371900 508358 372060
rect 338796 371700 339592 371702
rect 338796 371610 339791 371700
rect 150094 371535 150104 371595
rect 150164 371535 150189 371595
rect 150094 371525 150189 371535
rect 59829 371335 59914 371340
rect 59829 371280 59839 371335
rect 59904 371280 59914 371335
rect 59829 371265 59914 371280
rect 149829 371335 149914 371340
rect 149829 371280 149839 371335
rect 149904 371280 149914 371335
rect 149829 371265 149914 371280
rect 59829 370350 59911 371265
rect 49654 368640 49663 369730
rect 50753 368640 51258 369730
rect 52348 368640 52354 369730
rect 59769 369630 59979 370350
rect 68312 369730 68318 370600
rect 69188 369730 69194 370600
rect 149829 370350 149911 371265
rect 239451 370999 239546 371604
rect 239451 370939 239461 370999
rect 239521 370939 239546 370999
rect 239451 370929 239546 370939
rect 323888 371556 323970 371574
rect 323888 371500 323896 371556
rect 323964 371500 323970 371556
rect 239186 370739 239271 370744
rect 239186 370684 239196 370739
rect 239261 370684 239271 370739
rect 239186 370669 239271 370684
rect 57478 369420 61438 369630
rect 57478 366940 57688 369420
rect 61228 366965 61438 369420
rect 68318 369300 69188 369730
rect 139654 368640 139663 369730
rect 140753 368640 141258 369730
rect 142348 368640 142354 369730
rect 149769 369630 149979 370350
rect 158312 369730 158318 370600
rect 159188 369730 159194 370600
rect 239186 369754 239268 370669
rect 323888 370326 323970 371500
rect 338796 371364 338860 371610
rect 339000 371364 339791 371610
rect 338796 371282 339791 371364
rect 339192 371278 339791 371282
rect 340213 371278 340222 371700
rect 417544 371668 417598 371794
rect 417746 371786 418162 371794
rect 417746 371684 417996 371786
rect 418146 371684 418162 371786
rect 417746 371668 418162 371684
rect 417544 371638 418162 371668
rect 422664 371786 422866 371814
rect 420000 371642 420086 371650
rect 420000 371586 420008 371642
rect 420076 371586 420086 371642
rect 420000 371270 420086 371586
rect 420000 371206 420012 371270
rect 420084 371206 420086 371270
rect 420000 371189 420086 371206
rect 422664 371638 422696 371786
rect 422844 371638 422866 371786
rect 422664 371408 422866 371638
rect 422664 371204 422700 371408
rect 422830 371204 422866 371408
rect 508158 371300 508358 371900
rect 510358 372060 510558 372080
rect 510358 371900 510378 372060
rect 510538 372040 510558 372060
rect 510538 372030 510638 372040
rect 510538 371930 511088 372030
rect 510538 371920 510638 371930
rect 510538 371900 510558 371920
rect 510358 371880 510558 371900
rect 510988 371910 511088 371930
rect 511638 371940 511838 371960
rect 511638 371910 511658 371940
rect 509401 371844 509573 371864
rect 509401 371784 509441 371844
rect 509535 371784 509573 371844
rect 510988 371810 511658 371910
rect 509401 371756 509573 371784
rect 511638 371780 511658 371810
rect 511818 371780 511838 371940
rect 511638 371760 511838 371780
rect 509437 371542 509539 371756
rect 509437 371484 509445 371542
rect 509531 371484 509539 371542
rect 509437 371478 509539 371484
rect 422664 371178 422866 371204
rect 507518 371260 508358 371300
rect 507518 371140 507558 371260
rect 507758 371140 508358 371260
rect 507518 371100 508358 371140
rect 509437 371318 509539 371322
rect 509437 371260 509445 371318
rect 509531 371260 509539 371318
rect 509437 371014 509539 371260
rect 509397 370990 509569 371014
rect 509397 370930 509439 370990
rect 509533 370930 509569 370990
rect 509397 370906 509569 370930
rect 330798 370326 331758 370328
rect 147478 369420 151438 369630
rect 68318 368421 69188 368430
rect 57038 365130 58073 366940
rect 57038 364385 57193 365130
rect 57873 364385 58073 365130
rect 60793 365130 61758 366965
rect 147478 366940 147688 369420
rect 151228 366965 151438 369420
rect 158318 369300 159188 369730
rect 158318 368421 159188 368430
rect 237088 368517 238038 368525
rect 239126 368517 239336 369754
rect 247585 368633 247591 370134
rect 249092 368633 249098 370134
rect 323880 369374 331774 370326
rect 240798 368517 241743 368547
rect 237088 368178 241743 368517
rect 237088 368000 238038 368178
rect 60793 364385 60963 365130
rect 61643 364385 61758 365130
rect 147038 365130 148073 366940
rect 147038 364385 147193 365130
rect 147873 364385 148073 365130
rect 150793 365130 151758 366965
rect 150793 364385 150963 365130
rect 151643 364385 151758 365130
rect 237078 365900 238038 368000
rect 237078 365240 237258 365900
rect 237918 365240 238038 365900
rect 237078 365120 238038 365240
rect 240798 367812 241743 368178
rect 247591 368088 249092 368633
rect 240798 365900 241758 367812
rect 247591 366578 249092 366587
rect 240798 365240 240978 365900
rect 241638 365240 241758 365900
rect 240798 365120 241758 365240
rect 327078 365900 328038 369374
rect 327078 365240 327258 365900
rect 327918 365240 328038 365900
rect 327078 365120 328038 365240
rect 330798 365900 331758 369374
rect 330798 365240 330978 365900
rect 331638 365240 331758 365900
rect 330798 365120 331758 365240
rect 417078 368220 417238 368820
rect 417838 368220 418038 368820
rect 417078 365900 418038 368220
rect 417078 365240 417258 365900
rect 417918 365240 418038 365900
rect 417078 365120 418038 365240
rect 420798 368220 420958 368820
rect 421558 368220 421758 368820
rect 420798 365900 421758 368220
rect 420798 365240 420978 365900
rect 421638 365240 421758 365900
rect 420798 365120 421758 365240
rect 507078 368220 507238 368820
rect 507838 368220 508038 368820
rect 507078 365900 508038 368220
rect 507078 365240 507258 365900
rect 507918 365240 508038 365900
rect 507078 365120 508038 365240
rect 510798 368220 510958 368820
rect 511558 368220 511758 368820
rect 510798 365900 511758 368220
rect 510798 365240 510978 365900
rect 511638 365240 511758 365900
rect 510798 365120 511758 365240
rect 57038 364275 58073 364385
rect 147038 364275 148073 364385
rect 52344 360230 53664 360398
rect 52344 359406 52640 360230
rect 53366 359406 53664 360230
rect 52344 357788 53664 359406
rect 52344 357062 52608 357788
rect 53300 357062 53664 357788
rect 52344 356766 53664 357062
rect 142344 360230 143664 360398
rect 142344 359406 142640 360230
rect 143366 359406 143664 360230
rect 142344 357788 143664 359406
rect 142344 357062 142608 357788
rect 143300 357062 143664 357788
rect 142344 356766 143664 357062
rect 232344 360230 233664 360398
rect 232344 359406 232640 360230
rect 233366 359406 233664 360230
rect 232344 357788 233664 359406
rect 232344 357062 232608 357788
rect 233300 357062 233664 357788
rect 232344 356766 233664 357062
rect 322344 360230 323664 360398
rect 322344 359406 322640 360230
rect 323366 359406 323664 360230
rect 322344 357788 323664 359406
rect 322344 357062 322608 357788
rect 323300 357062 323664 357788
rect 322344 356766 323664 357062
rect 412344 360230 413664 360398
rect 412344 359406 412640 360230
rect 413366 359406 413664 360230
rect 412344 357788 413664 359406
rect 412344 357062 412608 357788
rect 413300 357062 413664 357788
rect 412344 356766 413664 357062
rect 502344 360230 503664 360398
rect 502344 359406 502640 360230
rect 503366 359406 503664 360230
rect 502344 357788 503664 359406
rect 502344 357062 502608 357788
rect 503300 357062 503664 357788
rect 502344 356766 503664 357062
rect 64428 266810 65748 267240
rect 64428 266084 64790 266810
rect 65482 266084 65748 266810
rect 64428 264794 65748 266084
rect 64428 263970 64790 264794
rect 65516 263970 65748 264794
rect 64428 263608 65748 263970
rect 153552 266606 154872 267036
rect 153552 265880 153914 266606
rect 154606 265880 154872 266606
rect 153552 264590 154872 265880
rect 153552 263766 153914 264590
rect 154640 263766 154872 264590
rect 153552 263404 154872 263766
rect 244806 266418 246126 266848
rect 244806 265692 245168 266418
rect 245860 265692 246126 266418
rect 244806 264402 246126 265692
rect 244806 263578 245168 264402
rect 245894 263578 246126 264402
rect 334428 266810 335748 267240
rect 334428 266084 334790 266810
rect 335482 266084 335748 266810
rect 334428 264794 335748 266084
rect 334428 263970 334790 264794
rect 335516 263970 335748 264794
rect 334428 263608 335748 263970
rect 424428 266810 425748 267240
rect 424428 266084 424790 266810
rect 425482 266084 425748 266810
rect 424428 264794 425748 266084
rect 424428 263970 424790 264794
rect 425516 263970 425748 264794
rect 424428 263608 425748 263970
rect 514428 266810 515748 267240
rect 514428 266084 514790 266810
rect 515482 266084 515748 266810
rect 514428 264794 515748 266084
rect 514428 263970 514790 264794
rect 515516 263970 515748 264794
rect 514428 263608 515748 263970
rect 244806 263216 246126 263578
rect 417108 259935 418093 260105
rect 417108 259190 417278 259935
rect 417958 259190 418093 259935
rect 417108 258510 418093 259190
rect 420828 259965 421828 260055
rect 420828 259220 420998 259965
rect 421678 259220 421828 259965
rect 57138 258380 58098 258500
rect 57138 257720 57318 258380
rect 57978 257720 58098 258380
rect 57138 255400 58098 257720
rect 57138 254800 57298 255400
rect 57898 254800 58098 255400
rect 60858 258380 61818 258500
rect 60858 257720 61038 258380
rect 61698 257720 61818 258380
rect 327138 258380 328098 258500
rect 60858 255400 61818 257720
rect 60858 254800 61018 255400
rect 61618 254800 61818 255400
rect 146262 258176 147222 258296
rect 146262 257516 146442 258176
rect 147102 257516 147222 258176
rect 146262 255196 147222 257516
rect 146262 254596 146422 255196
rect 147022 254596 147222 255196
rect 149982 258176 150942 258296
rect 149982 257516 150162 258176
rect 150822 257516 150942 258176
rect 149982 255196 150942 257516
rect 237516 257988 238476 258108
rect 237516 257328 237696 257988
rect 238356 257328 238476 257988
rect 237516 256437 238476 257328
rect 241236 257988 242196 258108
rect 241236 257328 241416 257988
rect 242076 257328 242196 257988
rect 241236 256437 242196 257328
rect 327138 257720 327318 258380
rect 327978 257720 328098 258380
rect 235106 256422 242205 256437
rect 149982 254596 150142 255196
rect 150742 254596 150942 255196
rect 234112 255365 242205 256422
rect 327138 255843 328098 257720
rect 330858 258380 331818 258500
rect 330858 257720 331038 258380
rect 331698 257720 331818 258380
rect 330858 255843 331818 257720
rect 417433 256895 417633 258510
rect 420828 258460 421828 259220
rect 507108 259935 508093 260105
rect 507108 259190 507278 259935
rect 507958 259190 508093 259935
rect 507108 258510 508093 259190
rect 510828 259965 511828 260055
rect 510828 259220 510998 259965
rect 511678 259220 511828 259965
rect 421203 256895 421403 258460
rect 417433 256695 421403 256895
rect 507433 256895 507633 258510
rect 510828 258460 511828 259220
rect 511203 256895 511403 258460
rect 507433 256695 511403 256895
rect 234112 253204 234674 255365
rect 327086 255282 331819 255843
rect 327138 255278 328098 255282
rect 320424 253495 320433 254443
rect 321381 253495 321390 254443
rect 234122 253110 234658 253204
rect 234122 252986 234286 253110
rect 234394 252986 234658 253110
rect 234122 252824 234658 252986
rect 320433 252790 321381 253495
rect 149124 252188 149210 252197
rect 149124 252124 149132 252188
rect 149204 252124 149210 252188
rect 58158 252060 58358 252080
rect 58158 251900 58178 252060
rect 58338 251900 58358 252060
rect 58158 251300 58358 251900
rect 60358 252060 60558 252080
rect 60358 251900 60378 252060
rect 60538 252040 60558 252060
rect 60538 252030 60638 252040
rect 60538 251930 61088 252030
rect 60538 251920 60638 251930
rect 60538 251900 60558 251920
rect 60358 251880 60558 251900
rect 60988 251910 61088 251930
rect 61638 251940 61838 251960
rect 61638 251910 61658 251940
rect 59401 251844 59573 251864
rect 59401 251784 59441 251844
rect 59535 251784 59573 251844
rect 60988 251810 61658 251910
rect 59401 251756 59573 251784
rect 61638 251780 61658 251810
rect 61818 251780 61838 251940
rect 61638 251760 61838 251780
rect 59437 251542 59539 251756
rect 149124 251668 149210 252124
rect 232171 251962 232497 251968
rect 59437 251484 59445 251542
rect 59531 251484 59539 251542
rect 59437 251478 59539 251484
rect 146668 251590 147286 251626
rect 149124 251612 149132 251668
rect 149200 251612 149210 251668
rect 231332 251636 231341 251962
rect 231667 251636 232171 251962
rect 320427 251842 320433 252790
rect 321381 251842 321387 252790
rect 232171 251630 232497 251636
rect 149124 251604 149210 251612
rect 146668 251464 146722 251590
rect 146870 251582 147286 251590
rect 146870 251480 147120 251582
rect 147270 251480 147286 251582
rect 146870 251464 147286 251480
rect 146668 251434 147286 251464
rect 151788 251582 151990 251610
rect 329396 251604 329596 255282
rect 330858 255261 331818 255282
rect 420039 252200 420239 256695
rect 510039 252200 510239 256695
rect 149124 251438 149210 251446
rect 149124 251382 149132 251438
rect 149200 251382 149210 251438
rect 57518 251260 58358 251300
rect 57518 251140 57558 251260
rect 57758 251140 58358 251260
rect 57518 251100 58358 251140
rect 59437 251318 59539 251322
rect 59437 251260 59445 251318
rect 59531 251260 59539 251318
rect 59437 251014 59539 251260
rect 149124 251066 149210 251382
rect 59397 250990 59569 251014
rect 59397 250930 59439 250990
rect 59533 250930 59569 250990
rect 149124 251002 149136 251066
rect 149208 251002 149210 251066
rect 149124 250985 149210 251002
rect 151788 251434 151820 251582
rect 151968 251434 151990 251582
rect 151788 251204 151990 251434
rect 151788 251000 151824 251204
rect 151954 251000 151990 251204
rect 249174 251308 249970 251310
rect 249174 251218 250169 251308
rect 151788 250974 151990 251000
rect 234266 251164 234348 251182
rect 234266 251108 234274 251164
rect 234342 251108 234348 251164
rect 59397 250906 59569 250930
rect 234266 249934 234348 251108
rect 249174 250972 249238 251218
rect 249378 250972 250169 251218
rect 249174 250890 250169 250972
rect 249570 250886 250169 250890
rect 250591 250886 250600 251308
rect 329451 250999 329546 251604
rect 420094 251595 420189 252200
rect 420094 251535 420104 251595
rect 420164 251535 420189 251595
rect 420094 251525 420189 251535
rect 510094 251595 510189 252200
rect 510094 251535 510104 251595
rect 510164 251535 510189 251595
rect 510094 251525 510189 251535
rect 329451 250939 329461 250999
rect 329521 250939 329546 250999
rect 329451 250929 329546 250939
rect 419829 251335 419914 251340
rect 419829 251280 419839 251335
rect 419904 251280 419914 251335
rect 419829 251265 419914 251280
rect 509829 251335 509914 251340
rect 509829 251280 509839 251335
rect 509904 251280 509914 251335
rect 509829 251265 509914 251280
rect 329186 250739 329271 250744
rect 329186 250684 329196 250739
rect 329261 250684 329271 250739
rect 329186 250669 329271 250684
rect 241176 249934 242136 249936
rect 234258 248982 242152 249934
rect 329186 249754 329268 250669
rect 419829 250350 419911 251265
rect 57078 248220 57238 248820
rect 57838 248220 58038 248820
rect 57078 245900 58038 248220
rect 57078 245240 57258 245900
rect 57918 245240 58038 245900
rect 57078 245120 58038 245240
rect 60798 248220 60958 248820
rect 61558 248220 61758 248820
rect 60798 245900 61758 248220
rect 60798 245240 60978 245900
rect 61638 245240 61758 245900
rect 60798 245120 61758 245240
rect 146202 248016 146362 248616
rect 146962 248016 147162 248616
rect 146202 245696 147162 248016
rect 146202 245036 146382 245696
rect 147042 245036 147162 245696
rect 146202 244916 147162 245036
rect 149922 248016 150082 248616
rect 150682 248016 150882 248616
rect 149922 245696 150882 248016
rect 149922 245036 150102 245696
rect 150762 245036 150882 245696
rect 149922 244916 150882 245036
rect 237456 245508 238416 248982
rect 237456 244848 237636 245508
rect 238296 244848 238416 245508
rect 237456 244728 238416 244848
rect 241176 245508 242136 248982
rect 327088 248517 328038 248525
rect 329126 248517 329336 249754
rect 337585 248633 337591 250134
rect 339092 248633 339098 250134
rect 409654 248640 409663 249730
rect 410753 248640 411258 249730
rect 412348 248640 412354 249730
rect 419769 249630 419979 250350
rect 428312 249730 428318 250600
rect 429188 249730 429194 250600
rect 509829 250350 509911 251265
rect 417478 249420 421438 249630
rect 330798 248517 331743 248547
rect 327088 248178 331743 248517
rect 327088 248000 328038 248178
rect 241176 244848 241356 245508
rect 242016 244848 242136 245508
rect 327078 245900 328038 248000
rect 327078 245240 327258 245900
rect 327918 245240 328038 245900
rect 327078 245120 328038 245240
rect 330798 247812 331743 248178
rect 337591 248088 339092 248633
rect 330798 245900 331758 247812
rect 417478 246940 417688 249420
rect 421228 246965 421438 249420
rect 428318 249300 429188 249730
rect 499654 248640 499663 249730
rect 500753 248640 501258 249730
rect 502348 248640 502354 249730
rect 509769 249630 509979 250350
rect 518312 249730 518318 250600
rect 519188 249730 519194 250600
rect 507478 249420 511438 249630
rect 428318 248421 429188 248430
rect 337591 246578 339092 246587
rect 330798 245240 330978 245900
rect 331638 245240 331758 245900
rect 330798 245120 331758 245240
rect 417038 245130 418073 246940
rect 241176 244728 242136 244848
rect 417038 244385 417193 245130
rect 417873 244385 418073 245130
rect 420793 245130 421758 246965
rect 507478 246940 507688 249420
rect 511228 246965 511438 249420
rect 518318 249300 519188 249730
rect 518318 248421 519188 248430
rect 420793 244385 420963 245130
rect 421643 244385 421758 245130
rect 507038 245130 508073 246940
rect 507038 244385 507193 245130
rect 507873 244385 508073 245130
rect 510793 245130 511758 246965
rect 510793 244385 510963 245130
rect 511643 244385 511758 245130
rect 417038 244275 418073 244385
rect 507038 244275 508073 244385
rect 52344 240230 53664 240398
rect 52344 239406 52640 240230
rect 53366 239406 53664 240230
rect 322344 240230 323664 240398
rect 52344 237788 53664 239406
rect 52344 237062 52608 237788
rect 53300 237062 53664 237788
rect 52344 236766 53664 237062
rect 141468 240026 142788 240194
rect 141468 239202 141764 240026
rect 142490 239202 142788 240026
rect 141468 237584 142788 239202
rect 141468 236858 141732 237584
rect 142424 236858 142788 237584
rect 141468 236562 142788 236858
rect 232722 239838 234042 240006
rect 232722 239014 233018 239838
rect 233744 239014 234042 239838
rect 232722 237396 234042 239014
rect 232722 236670 232986 237396
rect 233678 236670 234042 237396
rect 322344 239406 322640 240230
rect 323366 239406 323664 240230
rect 322344 237788 323664 239406
rect 322344 237062 322608 237788
rect 323300 237062 323664 237788
rect 322344 236766 323664 237062
rect 412344 240230 413664 240398
rect 412344 239406 412640 240230
rect 413366 239406 413664 240230
rect 412344 237788 413664 239406
rect 412344 237062 412608 237788
rect 413300 237062 413664 237788
rect 412344 236766 413664 237062
rect 502344 240230 503664 240398
rect 502344 239406 502640 240230
rect 503366 239406 503664 240230
rect 502344 237788 503664 239406
rect 502344 237062 502608 237788
rect 503300 237062 503664 237788
rect 502344 236766 503664 237062
rect 232722 236374 234042 236670
rect 57138 152280 58098 152400
rect 57138 151620 57318 152280
rect 57978 151620 58098 152280
rect 57138 149300 58098 151620
rect 57138 148700 57298 149300
rect 57898 148700 58098 149300
rect 60858 152280 61818 152400
rect 60858 151620 61038 152280
rect 61698 151620 61818 152280
rect 60858 149300 61818 151620
rect 60858 148700 61018 149300
rect 61618 148700 61818 149300
rect 147138 152280 148098 152400
rect 147138 151620 147318 152280
rect 147978 151620 148098 152280
rect 147138 149300 148098 151620
rect 147138 148700 147298 149300
rect 147898 148700 148098 149300
rect 150858 152280 151818 152400
rect 150858 151620 151038 152280
rect 151698 151620 151818 152280
rect 150858 149300 151818 151620
rect 150858 148700 151018 149300
rect 151618 148700 151818 149300
rect 237138 152280 238098 152400
rect 237138 151620 237318 152280
rect 237978 151620 238098 152280
rect 237138 149300 238098 151620
rect 237138 148700 237298 149300
rect 237898 148700 238098 149300
rect 240858 152280 241818 152400
rect 240858 151620 241038 152280
rect 241698 151620 241818 152280
rect 240858 149300 241818 151620
rect 240858 148700 241018 149300
rect 241618 148700 241818 149300
rect 327138 152280 328098 152400
rect 327138 151620 327318 152280
rect 327978 151620 328098 152280
rect 327138 149300 328098 151620
rect 327138 148700 327298 149300
rect 327898 148700 328098 149300
rect 330858 152280 331818 152400
rect 330858 151620 331038 152280
rect 331698 151620 331818 152280
rect 330858 149300 331818 151620
rect 330858 148700 331018 149300
rect 331618 148700 331818 149300
rect 417138 152280 418098 152400
rect 417138 151620 417318 152280
rect 417978 151620 418098 152280
rect 417138 149300 418098 151620
rect 417138 148700 417298 149300
rect 417898 148700 418098 149300
rect 420858 152280 421818 152400
rect 420858 151620 421038 152280
rect 421698 151620 421818 152280
rect 420858 149300 421818 151620
rect 420858 148700 421018 149300
rect 421618 148700 421818 149300
rect 507138 152280 508098 152400
rect 507138 151620 507318 152280
rect 507978 151620 508098 152280
rect 507138 149300 508098 151620
rect 507138 148700 507298 149300
rect 507898 148700 508098 149300
rect 510858 152280 511818 152400
rect 510858 151620 511038 152280
rect 511698 151620 511818 152280
rect 510858 149300 511818 151620
rect 510858 148700 511018 149300
rect 511618 148700 511818 149300
rect 58158 145960 58358 145980
rect 58158 145800 58178 145960
rect 58338 145800 58358 145960
rect 58158 145200 58358 145800
rect 60358 145960 60558 145980
rect 60358 145800 60378 145960
rect 60538 145940 60558 145960
rect 148158 145960 148358 145980
rect 60538 145930 60638 145940
rect 60538 145830 61088 145930
rect 60538 145820 60638 145830
rect 60538 145800 60558 145820
rect 60358 145780 60558 145800
rect 60988 145810 61088 145830
rect 61638 145840 61838 145860
rect 61638 145810 61658 145840
rect 60988 145710 61658 145810
rect 61638 145680 61658 145710
rect 61818 145680 61838 145840
rect 61638 145660 61838 145680
rect 148158 145800 148178 145960
rect 148338 145800 148358 145960
rect 148158 145200 148358 145800
rect 150358 145960 150558 145980
rect 150358 145800 150378 145960
rect 150538 145940 150558 145960
rect 238158 145960 238358 145980
rect 150538 145930 150638 145940
rect 150538 145830 151088 145930
rect 150538 145820 150638 145830
rect 150538 145800 150558 145820
rect 150358 145780 150558 145800
rect 150988 145810 151088 145830
rect 151638 145840 151838 145860
rect 151638 145810 151658 145840
rect 150988 145710 151658 145810
rect 151638 145680 151658 145710
rect 151818 145680 151838 145840
rect 151638 145660 151838 145680
rect 238158 145800 238178 145960
rect 238338 145800 238358 145960
rect 238158 145200 238358 145800
rect 240358 145960 240558 145980
rect 240358 145800 240378 145960
rect 240538 145940 240558 145960
rect 328158 145960 328358 145980
rect 240538 145930 240638 145940
rect 240538 145830 241088 145930
rect 240538 145820 240638 145830
rect 240538 145800 240558 145820
rect 240358 145780 240558 145800
rect 240988 145810 241088 145830
rect 241638 145840 241838 145860
rect 241638 145810 241658 145840
rect 240988 145710 241658 145810
rect 241638 145680 241658 145710
rect 241818 145680 241838 145840
rect 241638 145660 241838 145680
rect 328158 145800 328178 145960
rect 328338 145800 328358 145960
rect 328158 145200 328358 145800
rect 330358 145960 330558 145980
rect 330358 145800 330378 145960
rect 330538 145940 330558 145960
rect 418158 145960 418358 145980
rect 330538 145930 330638 145940
rect 330538 145830 331088 145930
rect 330538 145820 330638 145830
rect 330538 145800 330558 145820
rect 330358 145780 330558 145800
rect 330988 145810 331088 145830
rect 331638 145840 331838 145860
rect 331638 145810 331658 145840
rect 330988 145710 331658 145810
rect 331638 145680 331658 145710
rect 331818 145680 331838 145840
rect 331638 145660 331838 145680
rect 418158 145800 418178 145960
rect 418338 145800 418358 145960
rect 418158 145200 418358 145800
rect 420358 145960 420558 145980
rect 420358 145800 420378 145960
rect 420538 145940 420558 145960
rect 508158 145960 508358 145980
rect 420538 145930 420638 145940
rect 420538 145830 421088 145930
rect 420538 145820 420638 145830
rect 420538 145800 420558 145820
rect 420358 145780 420558 145800
rect 420988 145810 421088 145830
rect 421638 145840 421838 145860
rect 421638 145810 421658 145840
rect 420988 145710 421658 145810
rect 421638 145680 421658 145710
rect 421818 145680 421838 145840
rect 421638 145660 421838 145680
rect 508158 145800 508178 145960
rect 508338 145800 508358 145960
rect 508158 145200 508358 145800
rect 510358 145960 510558 145980
rect 510358 145800 510378 145960
rect 510538 145940 510558 145960
rect 510538 145930 510638 145940
rect 510538 145830 511088 145930
rect 510538 145820 510638 145830
rect 510538 145800 510558 145820
rect 510358 145780 510558 145800
rect 510988 145810 511088 145830
rect 511638 145840 511838 145860
rect 511638 145810 511658 145840
rect 510988 145710 511658 145810
rect 511638 145680 511658 145710
rect 511818 145680 511838 145840
rect 511638 145660 511838 145680
rect 57518 145160 58358 145200
rect 57518 145040 57558 145160
rect 57758 145040 58358 145160
rect 57518 145000 58358 145040
rect 147518 145160 148358 145200
rect 147518 145040 147558 145160
rect 147758 145040 148358 145160
rect 147518 145000 148358 145040
rect 237518 145160 238358 145200
rect 237518 145040 237558 145160
rect 237758 145040 238358 145160
rect 237518 145000 238358 145040
rect 327518 145160 328358 145200
rect 327518 145040 327558 145160
rect 327758 145040 328358 145160
rect 327518 145000 328358 145040
rect 417518 145160 418358 145200
rect 417518 145040 417558 145160
rect 417758 145040 418358 145160
rect 417518 145000 418358 145040
rect 507518 145160 508358 145200
rect 507518 145040 507558 145160
rect 507758 145040 508358 145160
rect 507518 145000 508358 145040
rect 57078 142120 57238 142720
rect 57838 142120 58038 142720
rect 57078 139800 58038 142120
rect 57078 139140 57258 139800
rect 57918 139140 58038 139800
rect 57078 139020 58038 139140
rect 60798 142120 60958 142720
rect 61558 142120 61758 142720
rect 60798 139800 61758 142120
rect 60798 139140 60978 139800
rect 61638 139140 61758 139800
rect 60798 139020 61758 139140
rect 147078 142120 147238 142720
rect 147838 142120 148038 142720
rect 147078 139800 148038 142120
rect 147078 139140 147258 139800
rect 147918 139140 148038 139800
rect 147078 139020 148038 139140
rect 150798 142120 150958 142720
rect 151558 142120 151758 142720
rect 150798 139800 151758 142120
rect 150798 139140 150978 139800
rect 151638 139140 151758 139800
rect 150798 139020 151758 139140
rect 237078 142120 237238 142720
rect 237838 142120 238038 142720
rect 237078 139800 238038 142120
rect 237078 139140 237258 139800
rect 237918 139140 238038 139800
rect 237078 139020 238038 139140
rect 240798 142120 240958 142720
rect 241558 142120 241758 142720
rect 240798 139800 241758 142120
rect 240798 139140 240978 139800
rect 241638 139140 241758 139800
rect 240798 139020 241758 139140
rect 327078 142120 327238 142720
rect 327838 142120 328038 142720
rect 327078 139800 328038 142120
rect 327078 139140 327258 139800
rect 327918 139140 328038 139800
rect 327078 139020 328038 139140
rect 330798 142120 330958 142720
rect 331558 142120 331758 142720
rect 330798 139800 331758 142120
rect 330798 139140 330978 139800
rect 331638 139140 331758 139800
rect 330798 139020 331758 139140
rect 417078 142120 417238 142720
rect 417838 142120 418038 142720
rect 417078 139800 418038 142120
rect 417078 139140 417258 139800
rect 417918 139140 418038 139800
rect 417078 139020 418038 139140
rect 420798 142120 420958 142720
rect 421558 142120 421758 142720
rect 420798 139800 421758 142120
rect 420798 139140 420978 139800
rect 421638 139140 421758 139800
rect 420798 139020 421758 139140
rect 507078 142120 507238 142720
rect 507838 142120 508038 142720
rect 507078 139800 508038 142120
rect 507078 139140 507258 139800
rect 507918 139140 508038 139800
rect 507078 139020 508038 139140
rect 510798 142120 510958 142720
rect 511558 142120 511758 142720
rect 510798 139800 511758 142120
rect 510798 139140 510978 139800
rect 511638 139140 511758 139800
rect 510798 139020 511758 139140
rect 57138 62280 58098 62400
rect 57138 61620 57318 62280
rect 57978 61620 58098 62280
rect 57138 59300 58098 61620
rect 57138 58700 57298 59300
rect 57898 58700 58098 59300
rect 60858 62280 61818 62400
rect 60858 61620 61038 62280
rect 61698 61620 61818 62280
rect 60858 59300 61818 61620
rect 60858 58700 61018 59300
rect 61618 58700 61818 59300
rect 147138 62280 148098 62400
rect 147138 61620 147318 62280
rect 147978 61620 148098 62280
rect 147138 59300 148098 61620
rect 147138 58700 147298 59300
rect 147898 58700 148098 59300
rect 150858 62280 151818 62400
rect 150858 61620 151038 62280
rect 151698 61620 151818 62280
rect 150858 59300 151818 61620
rect 150858 58700 151018 59300
rect 151618 58700 151818 59300
rect 237138 62280 238098 62400
rect 237138 61620 237318 62280
rect 237978 61620 238098 62280
rect 237138 59300 238098 61620
rect 237138 58700 237298 59300
rect 237898 58700 238098 59300
rect 240858 62280 241818 62400
rect 240858 61620 241038 62280
rect 241698 61620 241818 62280
rect 240858 59300 241818 61620
rect 240858 58700 241018 59300
rect 241618 58700 241818 59300
rect 327138 62280 328098 62400
rect 327138 61620 327318 62280
rect 327978 61620 328098 62280
rect 327138 59300 328098 61620
rect 327138 58700 327298 59300
rect 327898 58700 328098 59300
rect 330858 62280 331818 62400
rect 330858 61620 331038 62280
rect 331698 61620 331818 62280
rect 330858 59300 331818 61620
rect 330858 58700 331018 59300
rect 331618 58700 331818 59300
rect 417138 62280 418098 62400
rect 417138 61620 417318 62280
rect 417978 61620 418098 62280
rect 417138 59300 418098 61620
rect 417138 58700 417298 59300
rect 417898 58700 418098 59300
rect 420858 62280 421818 62400
rect 420858 61620 421038 62280
rect 421698 61620 421818 62280
rect 420858 59300 421818 61620
rect 420858 58700 421018 59300
rect 421618 58700 421818 59300
rect 507138 62280 508098 62400
rect 507138 61620 507318 62280
rect 507978 61620 508098 62280
rect 507138 59300 508098 61620
rect 507138 58700 507298 59300
rect 507898 58700 508098 59300
rect 510858 62280 511818 62400
rect 510858 61620 511038 62280
rect 511698 61620 511818 62280
rect 510858 59300 511818 61620
rect 510858 58700 511018 59300
rect 511618 58700 511818 59300
rect 58158 55960 58358 55980
rect 58158 55800 58178 55960
rect 58338 55800 58358 55960
rect 58158 55200 58358 55800
rect 60358 55960 60558 55980
rect 60358 55800 60378 55960
rect 60538 55940 60558 55960
rect 148158 55960 148358 55980
rect 60538 55930 60638 55940
rect 60538 55830 61088 55930
rect 60538 55820 60638 55830
rect 60538 55800 60558 55820
rect 60358 55780 60558 55800
rect 60988 55810 61088 55830
rect 61638 55840 61838 55860
rect 61638 55810 61658 55840
rect 60988 55710 61658 55810
rect 61638 55680 61658 55710
rect 61818 55680 61838 55840
rect 61638 55660 61838 55680
rect 148158 55800 148178 55960
rect 148338 55800 148358 55960
rect 148158 55200 148358 55800
rect 150358 55960 150558 55980
rect 150358 55800 150378 55960
rect 150538 55940 150558 55960
rect 238158 55960 238358 55980
rect 150538 55930 150638 55940
rect 150538 55830 151088 55930
rect 150538 55820 150638 55830
rect 150538 55800 150558 55820
rect 150358 55780 150558 55800
rect 150988 55810 151088 55830
rect 151638 55840 151838 55860
rect 151638 55810 151658 55840
rect 150988 55710 151658 55810
rect 151638 55680 151658 55710
rect 151818 55680 151838 55840
rect 151638 55660 151838 55680
rect 238158 55800 238178 55960
rect 238338 55800 238358 55960
rect 238158 55200 238358 55800
rect 240358 55960 240558 55980
rect 240358 55800 240378 55960
rect 240538 55940 240558 55960
rect 328158 55960 328358 55980
rect 240538 55930 240638 55940
rect 240538 55830 241088 55930
rect 240538 55820 240638 55830
rect 240538 55800 240558 55820
rect 240358 55780 240558 55800
rect 240988 55810 241088 55830
rect 241638 55840 241838 55860
rect 241638 55810 241658 55840
rect 240988 55710 241658 55810
rect 241638 55680 241658 55710
rect 241818 55680 241838 55840
rect 241638 55660 241838 55680
rect 328158 55800 328178 55960
rect 328338 55800 328358 55960
rect 328158 55200 328358 55800
rect 330358 55960 330558 55980
rect 330358 55800 330378 55960
rect 330538 55940 330558 55960
rect 418158 55960 418358 55980
rect 330538 55930 330638 55940
rect 330538 55830 331088 55930
rect 330538 55820 330638 55830
rect 330538 55800 330558 55820
rect 330358 55780 330558 55800
rect 330988 55810 331088 55830
rect 331638 55840 331838 55860
rect 331638 55810 331658 55840
rect 330988 55710 331658 55810
rect 331638 55680 331658 55710
rect 331818 55680 331838 55840
rect 331638 55660 331838 55680
rect 418158 55800 418178 55960
rect 418338 55800 418358 55960
rect 418158 55200 418358 55800
rect 420358 55960 420558 55980
rect 420358 55800 420378 55960
rect 420538 55940 420558 55960
rect 508158 55960 508358 55980
rect 420538 55930 420638 55940
rect 420538 55830 421088 55930
rect 420538 55820 420638 55830
rect 420538 55800 420558 55820
rect 420358 55780 420558 55800
rect 420988 55810 421088 55830
rect 421638 55840 421838 55860
rect 421638 55810 421658 55840
rect 420988 55710 421658 55810
rect 421638 55680 421658 55710
rect 421818 55680 421838 55840
rect 421638 55660 421838 55680
rect 508158 55800 508178 55960
rect 508338 55800 508358 55960
rect 508158 55200 508358 55800
rect 510358 55960 510558 55980
rect 510358 55800 510378 55960
rect 510538 55940 510558 55960
rect 510538 55930 510638 55940
rect 510538 55830 511088 55930
rect 510538 55820 510638 55830
rect 510538 55800 510558 55820
rect 510358 55780 510558 55800
rect 510988 55810 511088 55830
rect 511638 55840 511838 55860
rect 511638 55810 511658 55840
rect 510988 55710 511658 55810
rect 511638 55680 511658 55710
rect 511818 55680 511838 55840
rect 511638 55660 511838 55680
rect 57518 55160 58358 55200
rect 57518 55040 57558 55160
rect 57758 55040 58358 55160
rect 57518 55000 58358 55040
rect 147518 55160 148358 55200
rect 147518 55040 147558 55160
rect 147758 55040 148358 55160
rect 147518 55000 148358 55040
rect 237518 55160 238358 55200
rect 237518 55040 237558 55160
rect 237758 55040 238358 55160
rect 237518 55000 238358 55040
rect 327518 55160 328358 55200
rect 327518 55040 327558 55160
rect 327758 55040 328358 55160
rect 327518 55000 328358 55040
rect 417518 55160 418358 55200
rect 417518 55040 417558 55160
rect 417758 55040 418358 55160
rect 417518 55000 418358 55040
rect 507518 55160 508358 55200
rect 507518 55040 507558 55160
rect 507758 55040 508358 55160
rect 507518 55000 508358 55040
rect 57078 52120 57238 52720
rect 57838 52120 58038 52720
rect 57078 49800 58038 52120
rect 57078 49140 57258 49800
rect 57918 49140 58038 49800
rect 57078 49020 58038 49140
rect 60798 52120 60958 52720
rect 61558 52120 61758 52720
rect 60798 49800 61758 52120
rect 60798 49140 60978 49800
rect 61638 49140 61758 49800
rect 60798 49020 61758 49140
rect 147078 52120 147238 52720
rect 147838 52120 148038 52720
rect 147078 49800 148038 52120
rect 147078 49140 147258 49800
rect 147918 49140 148038 49800
rect 147078 49020 148038 49140
rect 150798 52120 150958 52720
rect 151558 52120 151758 52720
rect 150798 49800 151758 52120
rect 150798 49140 150978 49800
rect 151638 49140 151758 49800
rect 150798 49020 151758 49140
rect 237078 52120 237238 52720
rect 237838 52120 238038 52720
rect 237078 49800 238038 52120
rect 237078 49140 237258 49800
rect 237918 49140 238038 49800
rect 237078 49020 238038 49140
rect 240798 52120 240958 52720
rect 241558 52120 241758 52720
rect 240798 49800 241758 52120
rect 240798 49140 240978 49800
rect 241638 49140 241758 49800
rect 240798 49020 241758 49140
rect 327078 52120 327238 52720
rect 327838 52120 328038 52720
rect 327078 49800 328038 52120
rect 327078 49140 327258 49800
rect 327918 49140 328038 49800
rect 327078 49020 328038 49140
rect 330798 52120 330958 52720
rect 331558 52120 331758 52720
rect 330798 49800 331758 52120
rect 330798 49140 330978 49800
rect 331638 49140 331758 49800
rect 330798 49020 331758 49140
rect 417078 52120 417238 52720
rect 417838 52120 418038 52720
rect 417078 49800 418038 52120
rect 417078 49140 417258 49800
rect 417918 49140 418038 49800
rect 417078 49020 418038 49140
rect 420798 52120 420958 52720
rect 421558 52120 421758 52720
rect 420798 49800 421758 52120
rect 420798 49140 420978 49800
rect 421638 49140 421758 49800
rect 420798 49020 421758 49140
rect 507078 52120 507238 52720
rect 507838 52120 508038 52720
rect 507078 49800 508038 52120
rect 507078 49140 507258 49800
rect 507918 49140 508038 49800
rect 507078 49020 508038 49140
rect 510798 52120 510958 52720
rect 511558 52120 511758 52720
rect 510798 49800 511758 52120
rect 510798 49140 510978 49800
rect 511638 49140 511758 49800
rect 510798 49020 511758 49140
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 327120 663544 327780 664204
rect 57318 661620 57978 662280
rect 61038 661620 61698 662280
rect 147318 661620 147978 662280
rect 151038 661620 151698 662280
rect 237318 661620 237978 662280
rect 241038 661620 241698 662280
rect 330840 663544 331500 664204
rect 417120 663544 417780 664204
rect 420840 663544 421500 664204
rect 507120 663544 507780 664204
rect 510840 663544 511500 664204
rect 331460 657604 331620 657764
rect 421460 657604 421620 657764
rect 511460 657604 511620 657764
rect 327360 656964 327560 657084
rect 417360 656964 417560 657084
rect 507360 656964 507560 657084
rect 61658 655680 61818 655840
rect 151658 655680 151818 655840
rect 241658 655680 241818 655840
rect 57558 655040 57758 655160
rect 147558 655040 147758 655160
rect 237558 655040 237758 655160
rect 57258 649140 57918 649800
rect 60978 649140 61638 649800
rect 147258 649140 147918 649800
rect 150978 649140 151638 649800
rect 237258 649140 237918 649800
rect 327060 651064 327720 651724
rect 330780 651064 331440 651724
rect 417060 651064 417720 651724
rect 420780 651064 421440 651724
rect 507060 651064 507720 651724
rect 510780 651064 511440 651724
rect 240978 649140 241638 649800
rect 417120 588544 417780 589204
rect 57318 586620 57978 587280
rect 61038 586620 61698 587280
rect 147318 586620 147978 587280
rect 151038 586620 151698 587280
rect 237318 586620 237978 587280
rect 241038 586620 241698 587280
rect 327318 586620 327978 587280
rect 331038 586620 331698 587280
rect 420840 588544 421500 589204
rect 507120 588544 507780 589204
rect 510840 588544 511500 589204
rect 421460 582604 421620 582764
rect 511460 582604 511620 582764
rect 417360 581964 417560 582084
rect 507360 581964 507560 582084
rect 61658 580680 61818 580840
rect 151658 580680 151818 580840
rect 241658 580680 241818 580840
rect 331658 580680 331818 580840
rect 57558 580040 57758 580160
rect 147558 580040 147758 580160
rect 237558 580040 237758 580160
rect 327558 580040 327758 580160
rect 57258 574140 57918 574800
rect 60978 574140 61638 574800
rect 147258 574140 147918 574800
rect 150978 574140 151638 574800
rect 237258 574140 237918 574800
rect 240978 574140 241638 574800
rect 327258 574140 327918 574800
rect 417060 576064 417720 576724
rect 420780 576064 421440 576724
rect 507060 576064 507720 576724
rect 510780 576064 511440 576724
rect 330978 574140 331638 574800
rect 64790 506084 65482 506810
rect 154790 506084 155482 506810
rect 244790 506084 245482 506810
rect 334790 506084 335482 506810
rect 424790 506084 425482 506810
rect 514790 506084 515482 506810
rect 147278 499190 147958 499935
rect 150998 499220 151678 499965
rect 57318 497720 57978 498380
rect 61038 497720 61698 498380
rect 237318 497720 237978 498380
rect 241038 497720 241698 498380
rect 327318 497720 327978 498380
rect 331038 497720 331698 498380
rect 417318 497720 417978 498380
rect 230433 493495 231381 494443
rect 57598 491668 57746 491794
rect 421038 497720 421698 498380
rect 507318 497720 507978 498380
rect 511038 497720 511698 498380
rect 320963 492028 321289 492354
rect 62700 491204 62830 491408
rect 57258 485240 57918 485900
rect 139663 488640 140753 489730
rect 339791 491278 340213 491700
rect 421658 491780 421818 491940
rect 507598 491668 507746 491794
rect 417558 491140 417758 491260
rect 512700 491204 512830 491408
rect 158318 488430 159188 489300
rect 60978 485240 61638 485900
rect 147193 484385 147873 485130
rect 150963 484385 151643 485130
rect 237258 485240 237918 485900
rect 247591 486587 249092 488088
rect 240978 485240 241638 485900
rect 327258 485240 327918 485900
rect 330978 485240 331638 485900
rect 417258 485240 417918 485900
rect 420978 485240 421638 485900
rect 507258 485240 507918 485900
rect 510978 485240 511638 485900
rect 52608 477062 53300 477788
rect 142608 477062 143300 477788
rect 232608 477062 233300 477788
rect 322608 477062 323300 477788
rect 412608 477062 413300 477788
rect 502608 477062 503300 477788
rect 64790 386084 65482 386810
rect 154790 386084 155482 386810
rect 244790 386084 245482 386810
rect 334790 386084 335482 386810
rect 424790 386084 425482 386810
rect 514790 386084 515482 386810
rect 57278 379190 57958 379935
rect 60998 379220 61678 379965
rect 147278 379190 147958 379935
rect 150998 379220 151678 379965
rect 237318 377720 237978 378380
rect 241038 377720 241698 378380
rect 327318 377720 327978 378380
rect 331038 377720 331698 378380
rect 417318 377720 417978 378380
rect 230433 373495 231381 374443
rect 421038 377720 421698 378380
rect 507318 377720 507978 378380
rect 511038 377720 511698 378380
rect 320963 372028 321289 372354
rect 49663 368640 50753 369730
rect 68318 368430 69188 369300
rect 139663 368640 140753 369730
rect 339791 371278 340213 371700
rect 417598 371668 417746 371794
rect 422700 371204 422830 371408
rect 511658 371780 511818 371940
rect 507558 371140 507758 371260
rect 57193 364385 57873 365130
rect 158318 368430 159188 369300
rect 60963 364385 61643 365130
rect 147193 364385 147873 365130
rect 150963 364385 151643 365130
rect 237258 365240 237918 365900
rect 247591 366587 249092 368088
rect 240978 365240 241638 365900
rect 327258 365240 327918 365900
rect 330978 365240 331638 365900
rect 417258 365240 417918 365900
rect 420978 365240 421638 365900
rect 507258 365240 507918 365900
rect 510978 365240 511638 365900
rect 52608 357062 53300 357788
rect 142608 357062 143300 357788
rect 232608 357062 233300 357788
rect 322608 357062 323300 357788
rect 412608 357062 413300 357788
rect 502608 357062 503300 357788
rect 64790 266084 65482 266810
rect 153914 265880 154606 266606
rect 245168 265692 245860 266418
rect 334790 266084 335482 266810
rect 424790 266084 425482 266810
rect 514790 266084 515482 266810
rect 417278 259190 417958 259935
rect 420998 259220 421678 259965
rect 57318 257720 57978 258380
rect 61038 257720 61698 258380
rect 146442 257516 147102 258176
rect 150162 257516 150822 258176
rect 237696 257328 238356 257988
rect 241416 257328 242076 257988
rect 327318 257720 327978 258380
rect 331038 257720 331698 258380
rect 507278 259190 507958 259935
rect 510998 259220 511678 259965
rect 320433 253495 321381 254443
rect 61658 251780 61818 251940
rect 231341 251636 231667 251962
rect 146722 251464 146870 251590
rect 57558 251140 57758 251260
rect 151824 251000 151954 251204
rect 250169 250886 250591 251308
rect 57258 245240 57918 245900
rect 60978 245240 61638 245900
rect 146382 245036 147042 245696
rect 150102 245036 150762 245696
rect 237636 244848 238296 245508
rect 409663 248640 410753 249730
rect 241356 244848 242016 245508
rect 327258 245240 327918 245900
rect 337591 246587 339092 248088
rect 428318 248430 429188 249300
rect 499663 248640 500753 249730
rect 330978 245240 331638 245900
rect 417193 244385 417873 245130
rect 518318 248430 519188 249300
rect 420963 244385 421643 245130
rect 507193 244385 507873 245130
rect 510963 244385 511643 245130
rect 52608 237062 53300 237788
rect 141732 236858 142424 237584
rect 232986 236670 233678 237396
rect 322608 237062 323300 237788
rect 412608 237062 413300 237788
rect 502608 237062 503300 237788
rect 57318 151620 57978 152280
rect 61038 151620 61698 152280
rect 147318 151620 147978 152280
rect 151038 151620 151698 152280
rect 237318 151620 237978 152280
rect 241038 151620 241698 152280
rect 327318 151620 327978 152280
rect 331038 151620 331698 152280
rect 417318 151620 417978 152280
rect 421038 151620 421698 152280
rect 507318 151620 507978 152280
rect 511038 151620 511698 152280
rect 61658 145680 61818 145840
rect 151658 145680 151818 145840
rect 241658 145680 241818 145840
rect 331658 145680 331818 145840
rect 421658 145680 421818 145840
rect 511658 145680 511818 145840
rect 57558 145040 57758 145160
rect 147558 145040 147758 145160
rect 237558 145040 237758 145160
rect 327558 145040 327758 145160
rect 417558 145040 417758 145160
rect 507558 145040 507758 145160
rect 57258 139140 57918 139800
rect 60978 139140 61638 139800
rect 147258 139140 147918 139800
rect 150978 139140 151638 139800
rect 237258 139140 237918 139800
rect 240978 139140 241638 139800
rect 327258 139140 327918 139800
rect 330978 139140 331638 139800
rect 417258 139140 417918 139800
rect 420978 139140 421638 139800
rect 507258 139140 507918 139800
rect 510978 139140 511638 139800
rect 57318 61620 57978 62280
rect 61038 61620 61698 62280
rect 147318 61620 147978 62280
rect 151038 61620 151698 62280
rect 237318 61620 237978 62280
rect 241038 61620 241698 62280
rect 327318 61620 327978 62280
rect 331038 61620 331698 62280
rect 417318 61620 417978 62280
rect 421038 61620 421698 62280
rect 507318 61620 507978 62280
rect 511038 61620 511698 62280
rect 61658 55680 61818 55840
rect 151658 55680 151818 55840
rect 241658 55680 241818 55840
rect 331658 55680 331818 55840
rect 421658 55680 421818 55840
rect 511658 55680 511818 55840
rect 57558 55040 57758 55160
rect 147558 55040 147758 55160
rect 237558 55040 237758 55160
rect 327558 55040 327758 55160
rect 417558 55040 417758 55160
rect 507558 55040 507758 55160
rect 57258 49140 57918 49800
rect 60978 49140 61638 49800
rect 147258 49140 147918 49800
rect 150978 49140 151638 49800
rect 237258 49140 237918 49800
rect 240978 49140 241638 49800
rect 327258 49140 327918 49800
rect 330978 49140 331638 49800
rect 417258 49140 417918 49800
rect 420978 49140 421638 49800
rect 507258 49140 507918 49800
rect 510978 49140 511638 49800
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 702300 571594 704800
rect -800 680242 1700 685242
rect 582300 677984 584800 682984
rect 326940 667204 327900 667444
rect 326940 666424 327120 667204
rect 327780 666424 327900 667204
rect 57138 665280 58098 665520
rect 57138 664500 57318 665280
rect 57978 664500 58098 665280
rect 57138 662280 58098 664500
rect 57138 661620 57318 662280
rect 57978 661620 58098 662280
rect 57138 661440 58098 661620
rect 60858 665280 61818 665520
rect 60858 664500 61038 665280
rect 61698 664500 61818 665280
rect 60858 662280 61818 664500
rect 60858 661620 61038 662280
rect 61698 661620 61818 662280
rect 60858 661440 61818 661620
rect 147138 665280 148098 665520
rect 147138 664500 147318 665280
rect 147978 664500 148098 665280
rect 147138 662280 148098 664500
rect 147138 661620 147318 662280
rect 147978 661620 148098 662280
rect 147138 661440 148098 661620
rect 150858 665280 151818 665520
rect 150858 664500 151038 665280
rect 151698 664500 151818 665280
rect 150858 662280 151818 664500
rect 150858 661620 151038 662280
rect 151698 661620 151818 662280
rect 150858 661440 151818 661620
rect 237138 665280 238098 665520
rect 237138 664500 237318 665280
rect 237978 664500 238098 665280
rect 237138 662280 238098 664500
rect 237138 661620 237318 662280
rect 237978 661620 238098 662280
rect 237138 661440 238098 661620
rect 240858 665280 241818 665520
rect 240858 664500 241038 665280
rect 241698 664500 241818 665280
rect 240858 662280 241818 664500
rect 326940 664204 327900 666424
rect 326940 663544 327120 664204
rect 327780 663544 327900 664204
rect 326940 663364 327900 663544
rect 330660 667204 331620 667444
rect 330660 666424 330840 667204
rect 331500 666424 331620 667204
rect 330660 664204 331620 666424
rect 330660 663544 330840 664204
rect 331500 663544 331620 664204
rect 330660 663364 331620 663544
rect 416940 667204 417900 667444
rect 416940 666424 417120 667204
rect 417780 666424 417900 667204
rect 416940 664204 417900 666424
rect 416940 663544 417120 664204
rect 417780 663544 417900 664204
rect 416940 663364 417900 663544
rect 420660 667204 421620 667444
rect 420660 666424 420840 667204
rect 421500 666424 421620 667204
rect 420660 664204 421620 666424
rect 420660 663544 420840 664204
rect 421500 663544 421620 664204
rect 420660 663364 421620 663544
rect 506940 667204 507900 667444
rect 506940 666424 507120 667204
rect 507780 666424 507900 667204
rect 506940 664204 507900 666424
rect 506940 663544 507120 664204
rect 507780 663544 507900 664204
rect 506940 663364 507900 663544
rect 510660 667204 511620 667444
rect 510660 666424 510840 667204
rect 511500 666424 511620 667204
rect 510660 664204 511620 666424
rect 510660 663544 510840 664204
rect 511500 663544 511620 664204
rect 510660 663364 511620 663544
rect 240858 661620 241038 662280
rect 241698 661620 241818 662280
rect 240858 661440 241818 661620
rect 325636 657124 326868 657882
rect 331440 657764 331660 657784
rect 331440 657604 331460 657764
rect 331620 657762 331660 657764
rect 331620 657645 332777 657762
rect 333573 657645 334447 657665
rect 331620 657608 334447 657645
rect 331620 657604 331660 657608
rect 331440 657584 331660 657604
rect 332623 657364 334447 657608
rect 325636 656924 325686 657124
rect 325886 657084 327600 657124
rect 325886 656964 327360 657084
rect 327560 656964 327600 657084
rect 332623 657079 333750 657364
rect 325886 656924 327600 656964
rect 325636 656574 326868 656924
rect 332619 656914 333750 657079
rect 334200 656914 334447 657364
rect 332619 656629 334447 656914
rect 415636 657124 416868 657882
rect 421440 657764 421660 657784
rect 421440 657604 421460 657764
rect 421620 657762 421660 657764
rect 421620 657645 422777 657762
rect 423573 657645 424447 657665
rect 421620 657608 424447 657645
rect 421620 657604 421660 657608
rect 421440 657584 421660 657604
rect 422623 657364 424447 657608
rect 415636 656924 415686 657124
rect 415886 657084 417600 657124
rect 415886 656964 417360 657084
rect 417560 656964 417600 657084
rect 422623 657079 423750 657364
rect 415886 656924 417600 656964
rect 415636 656574 416868 656924
rect 422619 656914 423750 657079
rect 424200 656914 424447 657364
rect 422619 656629 424447 656914
rect 505636 657124 506868 657882
rect 511440 657764 511660 657784
rect 511440 657604 511460 657764
rect 511620 657762 511660 657764
rect 511620 657645 512777 657762
rect 513573 657645 514447 657665
rect 511620 657608 514447 657645
rect 511620 657604 511660 657608
rect 511440 657584 511660 657604
rect 512623 657364 514447 657608
rect 505636 656924 505686 657124
rect 505886 657084 507600 657124
rect 505886 656964 507360 657084
rect 507560 656964 507600 657084
rect 512623 657079 513750 657364
rect 505886 656924 507600 656964
rect 505636 656574 506868 656924
rect 512619 656914 513750 657079
rect 514200 656914 514447 657364
rect 512619 656629 514447 656914
rect 55834 655200 57066 655958
rect 61638 655840 61858 655860
rect 61638 655680 61658 655840
rect 61818 655838 61858 655840
rect 61818 655721 62975 655838
rect 63771 655721 64645 655741
rect 61818 655684 64645 655721
rect 61818 655680 61858 655684
rect 61638 655660 61858 655680
rect 62821 655440 64645 655684
rect 55834 655000 55884 655200
rect 56084 655160 57798 655200
rect 56084 655040 57558 655160
rect 57758 655040 57798 655160
rect 62821 655155 63948 655440
rect 56084 655000 57798 655040
rect 55834 654650 57066 655000
rect 62817 654990 63948 655155
rect 64398 654990 64645 655440
rect 62817 654705 64645 654990
rect 145834 655200 147066 655958
rect 151638 655840 151858 655860
rect 151638 655680 151658 655840
rect 151818 655838 151858 655840
rect 151818 655721 152975 655838
rect 153771 655721 154645 655741
rect 151818 655684 154645 655721
rect 151818 655680 151858 655684
rect 151638 655660 151858 655680
rect 152821 655440 154645 655684
rect 145834 655000 145884 655200
rect 146084 655160 147798 655200
rect 146084 655040 147558 655160
rect 147758 655040 147798 655160
rect 152821 655155 153948 655440
rect 146084 655000 147798 655040
rect 145834 654650 147066 655000
rect 152817 654990 153948 655155
rect 154398 654990 154645 655440
rect 152817 654705 154645 654990
rect 235834 655200 237066 655958
rect 241638 655840 241858 655860
rect 241638 655680 241658 655840
rect 241818 655838 241858 655840
rect 241818 655721 242975 655838
rect 243771 655721 244645 655741
rect 241818 655684 244645 655721
rect 241818 655680 241858 655684
rect 241638 655660 241858 655680
rect 242821 655440 244645 655684
rect 235834 655000 235884 655200
rect 236084 655160 237798 655200
rect 236084 655040 237558 655160
rect 237758 655040 237798 655160
rect 242821 655155 243948 655440
rect 236084 655000 237798 655040
rect 235834 654650 237066 655000
rect 242817 654990 243948 655155
rect 244398 654990 244645 655440
rect 242817 654705 244645 654990
rect 326880 651724 327840 651904
rect 326880 651064 327060 651724
rect 327720 651064 327840 651724
rect 57078 649800 58038 649980
rect 57078 649140 57258 649800
rect 57918 649140 58038 649800
rect -800 643842 1660 648642
rect 57078 646920 58038 649140
rect 57078 646140 57258 646920
rect 57918 646140 58038 646920
rect 57078 645900 58038 646140
rect 60798 649800 61758 649980
rect 60798 649140 60978 649800
rect 61638 649140 61758 649800
rect 60798 646920 61758 649140
rect 60798 646140 60978 646920
rect 61638 646140 61758 646920
rect 60798 645900 61758 646140
rect 147078 649800 148038 649980
rect 147078 649140 147258 649800
rect 147918 649140 148038 649800
rect 147078 646920 148038 649140
rect 147078 646140 147258 646920
rect 147918 646140 148038 646920
rect 147078 645900 148038 646140
rect 150798 649800 151758 649980
rect 150798 649140 150978 649800
rect 151638 649140 151758 649800
rect 150798 646920 151758 649140
rect 150798 646140 150978 646920
rect 151638 646140 151758 646920
rect 150798 645900 151758 646140
rect 237078 649800 238038 649980
rect 237078 649140 237258 649800
rect 237918 649140 238038 649800
rect 237078 646920 238038 649140
rect 237078 646140 237258 646920
rect 237918 646140 238038 646920
rect 237078 645900 238038 646140
rect 240798 649800 241758 649980
rect 240798 649140 240978 649800
rect 241638 649140 241758 649800
rect 240798 646920 241758 649140
rect 326880 648844 327840 651064
rect 326880 648064 327060 648844
rect 327720 648064 327840 648844
rect 326880 647824 327840 648064
rect 330600 651724 331560 651904
rect 330600 651064 330780 651724
rect 331440 651064 331560 651724
rect 330600 648844 331560 651064
rect 330600 648064 330780 648844
rect 331440 648064 331560 648844
rect 330600 647824 331560 648064
rect 416880 651724 417840 651904
rect 416880 651064 417060 651724
rect 417720 651064 417840 651724
rect 416880 648844 417840 651064
rect 416880 648064 417060 648844
rect 417720 648064 417840 648844
rect 416880 647824 417840 648064
rect 420600 651724 421560 651904
rect 420600 651064 420780 651724
rect 421440 651064 421560 651724
rect 420600 648844 421560 651064
rect 420600 648064 420780 648844
rect 421440 648064 421560 648844
rect 420600 647824 421560 648064
rect 506880 651724 507840 651904
rect 506880 651064 507060 651724
rect 507720 651064 507840 651724
rect 506880 648844 507840 651064
rect 506880 648064 507060 648844
rect 507720 648064 507840 648844
rect 506880 647824 507840 648064
rect 510600 651724 511560 651904
rect 510600 651064 510780 651724
rect 511440 651064 511560 651724
rect 510600 648844 511560 651064
rect 510600 648064 510780 648844
rect 511440 648064 511560 648844
rect 510600 647824 511560 648064
rect 240798 646140 240978 646920
rect 241638 646140 241758 646920
rect 240798 645900 241758 646140
rect 582340 639784 584800 644584
rect -800 633842 1660 638642
rect 582340 629784 584800 634584
rect 416940 592204 417900 592444
rect 416940 591424 417120 592204
rect 417780 591424 417900 592204
rect 57138 590280 58098 590520
rect 57138 589500 57318 590280
rect 57978 589500 58098 590280
rect 57138 587280 58098 589500
rect 57138 586620 57318 587280
rect 57978 586620 58098 587280
rect 57138 586440 58098 586620
rect 60858 590280 61818 590520
rect 60858 589500 61038 590280
rect 61698 589500 61818 590280
rect 60858 587280 61818 589500
rect 60858 586620 61038 587280
rect 61698 586620 61818 587280
rect 60858 586440 61818 586620
rect 147138 590280 148098 590520
rect 147138 589500 147318 590280
rect 147978 589500 148098 590280
rect 147138 587280 148098 589500
rect 147138 586620 147318 587280
rect 147978 586620 148098 587280
rect 147138 586440 148098 586620
rect 150858 590280 151818 590520
rect 150858 589500 151038 590280
rect 151698 589500 151818 590280
rect 150858 587280 151818 589500
rect 150858 586620 151038 587280
rect 151698 586620 151818 587280
rect 150858 586440 151818 586620
rect 237138 590280 238098 590520
rect 237138 589500 237318 590280
rect 237978 589500 238098 590280
rect 237138 587280 238098 589500
rect 237138 586620 237318 587280
rect 237978 586620 238098 587280
rect 237138 586440 238098 586620
rect 240858 590280 241818 590520
rect 240858 589500 241038 590280
rect 241698 589500 241818 590280
rect 240858 587280 241818 589500
rect 240858 586620 241038 587280
rect 241698 586620 241818 587280
rect 240858 586440 241818 586620
rect 327138 590280 328098 590520
rect 327138 589500 327318 590280
rect 327978 589500 328098 590280
rect 327138 587280 328098 589500
rect 327138 586620 327318 587280
rect 327978 586620 328098 587280
rect 327138 586440 328098 586620
rect 330858 590280 331818 590520
rect 330858 589500 331038 590280
rect 331698 589500 331818 590280
rect 330858 587280 331818 589500
rect 416940 589204 417900 591424
rect 416940 588544 417120 589204
rect 417780 588544 417900 589204
rect 416940 588364 417900 588544
rect 420660 592204 421620 592444
rect 420660 591424 420840 592204
rect 421500 591424 421620 592204
rect 420660 589204 421620 591424
rect 420660 588544 420840 589204
rect 421500 588544 421620 589204
rect 420660 588364 421620 588544
rect 506940 592204 507900 592444
rect 506940 591424 507120 592204
rect 507780 591424 507900 592204
rect 506940 589204 507900 591424
rect 506940 588544 507120 589204
rect 507780 588544 507900 589204
rect 506940 588364 507900 588544
rect 510660 592204 511620 592444
rect 510660 591424 510840 592204
rect 511500 591424 511620 592204
rect 510660 589204 511620 591424
rect 583520 589472 584800 589584
rect 510660 588544 510840 589204
rect 511500 588544 511620 589204
rect 510660 588364 511620 588544
rect 583520 588290 584800 588402
rect 330858 586620 331038 587280
rect 331698 586620 331818 587280
rect 583520 587108 584800 587220
rect 330858 586440 331818 586620
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 415636 582124 416868 582882
rect 421440 582764 421660 582784
rect 421440 582604 421460 582764
rect 421620 582762 421660 582764
rect 421620 582645 422777 582762
rect 423573 582645 424447 582665
rect 421620 582608 424447 582645
rect 421620 582604 421660 582608
rect 421440 582584 421660 582604
rect 422623 582364 424447 582608
rect 415636 581924 415686 582124
rect 415886 582084 417600 582124
rect 415886 581964 417360 582084
rect 417560 581964 417600 582084
rect 422623 582079 423750 582364
rect 415886 581924 417600 581964
rect 415636 581574 416868 581924
rect 422619 581914 423750 582079
rect 424200 581914 424447 582364
rect 422619 581629 424447 581914
rect 505636 582124 506868 582882
rect 511440 582764 511660 582784
rect 511440 582604 511460 582764
rect 511620 582762 511660 582764
rect 511620 582645 512777 582762
rect 513573 582645 514447 582665
rect 511620 582608 514447 582645
rect 511620 582604 511660 582608
rect 511440 582584 511660 582604
rect 512623 582364 514447 582608
rect 505636 581924 505686 582124
rect 505886 582084 507600 582124
rect 505886 581964 507360 582084
rect 507560 581964 507600 582084
rect 512623 582079 513750 582364
rect 505886 581924 507600 581964
rect 505636 581574 506868 581924
rect 512619 581914 513750 582079
rect 514200 581914 514447 582364
rect 512619 581629 514447 581914
rect 55834 580200 57066 580958
rect 61638 580840 61858 580860
rect 61638 580680 61658 580840
rect 61818 580838 61858 580840
rect 61818 580721 62975 580838
rect 63771 580721 64645 580741
rect 61818 580684 64645 580721
rect 61818 580680 61858 580684
rect 61638 580660 61858 580680
rect 62821 580440 64645 580684
rect 55834 580000 55884 580200
rect 56084 580160 57798 580200
rect 56084 580040 57558 580160
rect 57758 580040 57798 580160
rect 62821 580155 63948 580440
rect 56084 580000 57798 580040
rect 55834 579650 57066 580000
rect 62817 579990 63948 580155
rect 64398 579990 64645 580440
rect 62817 579705 64645 579990
rect 145834 580200 147066 580958
rect 151638 580840 151858 580860
rect 151638 580680 151658 580840
rect 151818 580838 151858 580840
rect 151818 580721 152975 580838
rect 153771 580721 154645 580741
rect 151818 580684 154645 580721
rect 151818 580680 151858 580684
rect 151638 580660 151858 580680
rect 152821 580440 154645 580684
rect 145834 580000 145884 580200
rect 146084 580160 147798 580200
rect 146084 580040 147558 580160
rect 147758 580040 147798 580160
rect 152821 580155 153948 580440
rect 146084 580000 147798 580040
rect 145834 579650 147066 580000
rect 152817 579990 153948 580155
rect 154398 579990 154645 580440
rect 152817 579705 154645 579990
rect 235834 580200 237066 580958
rect 241638 580840 241858 580860
rect 241638 580680 241658 580840
rect 241818 580838 241858 580840
rect 241818 580721 242975 580838
rect 243771 580721 244645 580741
rect 241818 580684 244645 580721
rect 241818 580680 241858 580684
rect 241638 580660 241858 580680
rect 242821 580440 244645 580684
rect 235834 580000 235884 580200
rect 236084 580160 237798 580200
rect 236084 580040 237558 580160
rect 237758 580040 237798 580160
rect 242821 580155 243948 580440
rect 236084 580000 237798 580040
rect 235834 579650 237066 580000
rect 242817 579990 243948 580155
rect 244398 579990 244645 580440
rect 242817 579705 244645 579990
rect 325834 580200 327066 580958
rect 331638 580840 331858 580860
rect 331638 580680 331658 580840
rect 331818 580838 331858 580840
rect 331818 580721 332975 580838
rect 333771 580721 334645 580741
rect 331818 580684 334645 580721
rect 331818 580680 331858 580684
rect 331638 580660 331858 580680
rect 332821 580440 334645 580684
rect 325834 580000 325884 580200
rect 326084 580160 327798 580200
rect 326084 580040 327558 580160
rect 327758 580040 327798 580160
rect 332821 580155 333948 580440
rect 326084 580000 327798 580040
rect 325834 579650 327066 580000
rect 332817 579990 333948 580155
rect 334398 579990 334645 580440
rect 332817 579705 334645 579990
rect 416880 576724 417840 576904
rect 416880 576064 417060 576724
rect 417720 576064 417840 576724
rect 57078 574800 58038 574980
rect 57078 574140 57258 574800
rect 57918 574140 58038 574800
rect 57078 571920 58038 574140
rect 57078 571140 57258 571920
rect 57918 571140 58038 571920
rect 57078 570900 58038 571140
rect 60798 574800 61758 574980
rect 60798 574140 60978 574800
rect 61638 574140 61758 574800
rect 60798 571920 61758 574140
rect 60798 571140 60978 571920
rect 61638 571140 61758 571920
rect 60798 570900 61758 571140
rect 147078 574800 148038 574980
rect 147078 574140 147258 574800
rect 147918 574140 148038 574800
rect 147078 571920 148038 574140
rect 147078 571140 147258 571920
rect 147918 571140 148038 571920
rect 147078 570900 148038 571140
rect 150798 574800 151758 574980
rect 150798 574140 150978 574800
rect 151638 574140 151758 574800
rect 150798 571920 151758 574140
rect 150798 571140 150978 571920
rect 151638 571140 151758 571920
rect 150798 570900 151758 571140
rect 237078 574800 238038 574980
rect 237078 574140 237258 574800
rect 237918 574140 238038 574800
rect 237078 571920 238038 574140
rect 237078 571140 237258 571920
rect 237918 571140 238038 571920
rect 237078 570900 238038 571140
rect 240798 574800 241758 574980
rect 240798 574140 240978 574800
rect 241638 574140 241758 574800
rect 240798 571920 241758 574140
rect 240798 571140 240978 571920
rect 241638 571140 241758 571920
rect 240798 570900 241758 571140
rect 327078 574800 328038 574980
rect 327078 574140 327258 574800
rect 327918 574140 328038 574800
rect 327078 571920 328038 574140
rect 327078 571140 327258 571920
rect 327918 571140 328038 571920
rect 327078 570900 328038 571140
rect 330798 574800 331758 574980
rect 330798 574140 330978 574800
rect 331638 574140 331758 574800
rect 330798 571920 331758 574140
rect 416880 573844 417840 576064
rect 416880 573064 417060 573844
rect 417720 573064 417840 573844
rect 416880 572824 417840 573064
rect 420600 576724 421560 576904
rect 420600 576064 420780 576724
rect 421440 576064 421560 576724
rect 420600 573844 421560 576064
rect 420600 573064 420780 573844
rect 421440 573064 421560 573844
rect 420600 572824 421560 573064
rect 506880 576724 507840 576904
rect 506880 576064 507060 576724
rect 507720 576064 507840 576724
rect 506880 573844 507840 576064
rect 506880 573064 507060 573844
rect 507720 573064 507840 573844
rect 506880 572824 507840 573064
rect 510600 576724 511560 576904
rect 510600 576064 510780 576724
rect 511440 576064 511560 576724
rect 510600 573844 511560 576064
rect 510600 573064 510780 573844
rect 511440 573064 511560 573844
rect 510600 572824 511560 573064
rect 330798 571140 330978 571920
rect 331638 571140 331758 571920
rect 330798 570900 331758 571140
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect -800 511530 480 511642
rect -800 510348 480 510460
rect 64524 509424 65714 509832
rect -800 509166 480 509278
rect 64524 508500 64750 509424
rect 65426 508500 65714 509424
rect -800 507984 480 508096
rect -800 506802 480 506914
rect 64524 506810 65714 508500
rect 64524 506084 64790 506810
rect 65482 506084 65714 506810
rect 64524 505736 65714 506084
rect 154524 509424 155714 509832
rect 154524 508500 154750 509424
rect 155426 508500 155714 509424
rect 154524 506810 155714 508500
rect 154524 506084 154790 506810
rect 155482 506084 155714 506810
rect 154524 505736 155714 506084
rect 244524 509424 245714 509832
rect 244524 508500 244750 509424
rect 245426 508500 245714 509424
rect 244524 506810 245714 508500
rect 244524 506084 244790 506810
rect 245482 506084 245714 506810
rect 244524 505736 245714 506084
rect 334524 509424 335714 509832
rect 334524 508500 334750 509424
rect 335426 508500 335714 509424
rect 334524 506810 335714 508500
rect 334524 506084 334790 506810
rect 335482 506084 335714 506810
rect 334524 505736 335714 506084
rect 424524 509424 425714 509832
rect 424524 508500 424750 509424
rect 425426 508500 425714 509424
rect 424524 506810 425714 508500
rect 424524 506084 424790 506810
rect 425482 506084 425714 506810
rect 424524 505736 425714 506084
rect 514524 509424 515714 509832
rect 514524 508500 514750 509424
rect 515426 508500 515714 509424
rect 514524 506810 515714 508500
rect 514524 506084 514790 506810
rect 515482 506084 515714 506810
rect 514524 505736 515714 506084
rect -800 505620 480 505732
rect 57138 501380 58098 501620
rect 57138 500600 57318 501380
rect 57978 500600 58098 501380
rect 57138 498380 58098 500600
rect 57138 497720 57318 498380
rect 57978 497720 58098 498380
rect 57138 497540 58098 497720
rect 60858 501380 61818 501620
rect 60858 500600 61038 501380
rect 61698 500600 61818 501380
rect 60858 498380 61818 500600
rect 147138 501380 148098 501620
rect 147138 500600 147318 501380
rect 147978 500600 148098 501380
rect 147138 499935 148098 500600
rect 147138 499190 147278 499935
rect 147958 499190 148098 499935
rect 147138 498735 148098 499190
rect 150858 501380 151818 501620
rect 150858 500600 151038 501380
rect 151698 500600 151818 501380
rect 150858 499965 151818 500600
rect 150858 499220 150998 499965
rect 151678 499220 151818 499965
rect 150858 498735 151818 499220
rect 237138 501380 238098 501620
rect 237138 500600 237318 501380
rect 237978 500600 238098 501380
rect 60858 497720 61038 498380
rect 61698 497720 61818 498380
rect 60858 497540 61818 497720
rect 237138 498380 238098 500600
rect 237138 497720 237318 498380
rect 237978 497720 238098 498380
rect 237138 497540 238098 497720
rect 240858 501380 241818 501620
rect 240858 500600 241038 501380
rect 241698 500600 241818 501380
rect 240858 498380 241818 500600
rect 240858 497720 241038 498380
rect 241698 497720 241818 498380
rect 240858 497540 241818 497720
rect 327138 501380 328098 501620
rect 327138 500600 327318 501380
rect 327978 500600 328098 501380
rect 327138 498380 328098 500600
rect 327138 497720 327318 498380
rect 327978 497720 328098 498380
rect 327138 497540 328098 497720
rect 330858 501380 331818 501620
rect 330858 500600 331038 501380
rect 331698 500600 331818 501380
rect 330858 498380 331818 500600
rect 330858 497720 331038 498380
rect 331698 497720 331818 498380
rect 330858 497540 331818 497720
rect 417138 501380 418098 501620
rect 417138 500600 417318 501380
rect 417978 500600 418098 501380
rect 417138 498380 418098 500600
rect 417138 497720 417318 498380
rect 417978 497720 418098 498380
rect 417138 497540 418098 497720
rect 420858 501380 421818 501620
rect 420858 500600 421038 501380
rect 421698 500600 421818 501380
rect 420858 498380 421818 500600
rect 420858 497720 421038 498380
rect 421698 497720 421818 498380
rect 420858 497540 421818 497720
rect 507138 501380 508098 501620
rect 507138 500600 507318 501380
rect 507978 500600 508098 501380
rect 507138 498380 508098 500600
rect 507138 497720 507318 498380
rect 507978 497720 508098 498380
rect 507138 497540 508098 497720
rect 510858 501380 511818 501620
rect 510858 500600 511038 501380
rect 511698 500600 511818 501380
rect 510858 498380 511818 500600
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 510858 497720 511038 498380
rect 511698 497720 511818 498380
rect 510858 497540 511818 497720
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 230428 494443 231386 494448
rect 229045 493495 229051 494443
rect 229999 493495 230433 494443
rect 231381 493495 231386 494443
rect 583520 494140 584800 494252
rect 230428 493490 231386 493495
rect 320958 492354 321294 492359
rect 55834 491300 57066 492058
rect 320269 492028 320275 492354
rect 320601 492028 320963 492354
rect 321289 492028 321294 492354
rect 320958 492023 321294 492028
rect 57542 491794 57798 491830
rect 63771 491821 64645 491841
rect 57542 491668 57598 491794
rect 57746 491668 57798 491794
rect 55834 491100 55884 491300
rect 56084 491294 57284 491300
rect 57542 491294 57798 491668
rect 63278 491540 64645 491821
rect 63278 491486 63948 491540
rect 56084 491100 57798 491294
rect 62664 491408 63948 491486
rect 62664 491204 62700 491408
rect 62830 491204 63948 491408
rect 62664 491172 63948 491204
rect 55834 490750 57066 491100
rect 57216 491094 57798 491100
rect 57542 491092 57798 491094
rect 63278 491090 63948 491172
rect 64398 491090 64645 491540
rect 339786 491700 340218 491705
rect 339786 491278 339791 491700
rect 340213 491278 340369 491700
rect 340791 491278 340797 491700
rect 415834 491300 417066 492058
rect 421638 491940 421858 491960
rect 421638 491780 421658 491940
rect 421818 491938 421858 491940
rect 421818 491821 422975 491938
rect 423771 491821 424645 491841
rect 421818 491784 424645 491821
rect 421818 491780 421858 491784
rect 421638 491760 421858 491780
rect 422821 491540 424645 491784
rect 339786 491273 340218 491278
rect 63278 490805 64645 491090
rect 415834 491100 415884 491300
rect 416084 491260 417798 491300
rect 416084 491140 417558 491260
rect 417758 491140 417798 491260
rect 422821 491255 423948 491540
rect 416084 491100 417798 491140
rect 415834 490750 417066 491100
rect 422817 491090 423948 491255
rect 424398 491090 424645 491540
rect 422817 490805 424645 491090
rect 505834 491300 507066 492058
rect 507542 491794 507798 491830
rect 513771 491821 514645 491841
rect 507542 491668 507598 491794
rect 507746 491668 507798 491794
rect 505834 491100 505884 491300
rect 506084 491294 507284 491300
rect 507542 491294 507798 491668
rect 513278 491540 514645 491821
rect 513278 491486 513948 491540
rect 506084 491100 507798 491294
rect 512664 491408 513948 491486
rect 512664 491204 512700 491408
rect 512830 491204 513948 491408
rect 512664 491172 513948 491204
rect 505834 490750 507066 491100
rect 507216 491094 507798 491100
rect 507542 491092 507798 491094
rect 513278 491090 513948 491172
rect 514398 491090 514645 491540
rect 513278 490805 514645 491090
rect 139658 489730 140758 489735
rect 139658 488640 139663 489730
rect 140753 488640 140758 489730
rect 139658 488635 140758 488640
rect 158313 489300 159193 489305
rect 139663 487805 140753 488635
rect 158313 488430 158318 489300
rect 159188 488430 159193 489300
rect 158313 488425 159193 488430
rect 139663 486709 140753 486715
rect 158318 487410 159188 488425
rect 247586 488089 249097 488093
rect 247586 488088 249825 488089
rect 247586 486587 247591 488088
rect 249092 486588 249825 488088
rect 251326 486588 251332 488089
rect 249092 486587 249097 486588
rect 247586 486582 249097 486587
rect 158318 486534 159188 486540
rect 57078 485900 58038 486080
rect 57078 485240 57258 485900
rect 57918 485240 58038 485900
rect 57078 483020 58038 485240
rect 57078 482240 57258 483020
rect 57918 482240 58038 483020
rect 57078 482000 58038 482240
rect 60798 485900 61758 486080
rect 60798 485240 60978 485900
rect 61638 485240 61758 485900
rect 237078 485900 238038 486080
rect 60798 483020 61758 485240
rect 147073 485130 148033 485275
rect 237078 485240 237258 485900
rect 237918 485240 238038 485900
rect 147073 484385 147193 485130
rect 147873 484665 148033 485130
rect 150798 485130 151758 485220
rect 147873 484385 148038 484665
rect 147073 484315 148038 484385
rect 60798 482240 60978 483020
rect 61638 482240 61758 483020
rect 60798 482000 61758 482240
rect 147078 483020 148038 484315
rect 147078 482240 147258 483020
rect 147918 482240 148038 483020
rect 147078 482000 148038 482240
rect 150798 484385 150963 485130
rect 151643 484385 151758 485130
rect 150798 483020 151758 484385
rect 150798 482240 150978 483020
rect 151638 482240 151758 483020
rect 150798 482000 151758 482240
rect 237078 483020 238038 485240
rect 237078 482240 237258 483020
rect 237918 482240 238038 483020
rect 237078 482000 238038 482240
rect 240798 485900 241758 486080
rect 240798 485240 240978 485900
rect 241638 485240 241758 485900
rect 240798 483020 241758 485240
rect 240798 482240 240978 483020
rect 241638 482240 241758 483020
rect 240798 482000 241758 482240
rect 327078 485900 328038 486080
rect 327078 485240 327258 485900
rect 327918 485240 328038 485900
rect 327078 483020 328038 485240
rect 327078 482240 327258 483020
rect 327918 482240 328038 483020
rect 327078 482000 328038 482240
rect 330798 485900 331758 486080
rect 330798 485240 330978 485900
rect 331638 485240 331758 485900
rect 330798 483020 331758 485240
rect 330798 482240 330978 483020
rect 331638 482240 331758 483020
rect 330798 482000 331758 482240
rect 417078 485900 418038 486080
rect 417078 485240 417258 485900
rect 417918 485240 418038 485900
rect 417078 483020 418038 485240
rect 417078 482240 417258 483020
rect 417918 482240 418038 483020
rect 417078 482000 418038 482240
rect 420798 485900 421758 486080
rect 420798 485240 420978 485900
rect 421638 485240 421758 485900
rect 420798 483020 421758 485240
rect 420798 482240 420978 483020
rect 421638 482240 421758 483020
rect 420798 482000 421758 482240
rect 507078 485900 508038 486080
rect 507078 485240 507258 485900
rect 507918 485240 508038 485900
rect 507078 483020 508038 485240
rect 507078 482240 507258 483020
rect 507918 482240 508038 483020
rect 507078 482000 508038 482240
rect 510798 485900 511758 486080
rect 510798 485240 510978 485900
rect 511638 485240 511758 485900
rect 510798 483020 511758 485240
rect 510798 482240 510978 483020
rect 511638 482240 511758 483020
rect 510798 482000 511758 482240
rect 52344 477788 53534 477990
rect 52344 477062 52608 477788
rect 53300 477062 53534 477788
rect 52344 475098 53534 477062
rect 52344 474174 52604 475098
rect 53280 474174 53534 475098
rect 52344 473894 53534 474174
rect 142344 477788 143534 477990
rect 142344 477062 142608 477788
rect 143300 477062 143534 477788
rect 142344 475098 143534 477062
rect 142344 474174 142604 475098
rect 143280 474174 143534 475098
rect 142344 473894 143534 474174
rect 232344 477788 233534 477990
rect 232344 477062 232608 477788
rect 233300 477062 233534 477788
rect 232344 475098 233534 477062
rect 232344 474174 232604 475098
rect 233280 474174 233534 475098
rect 232344 473894 233534 474174
rect 322344 477788 323534 477990
rect 322344 477062 322608 477788
rect 323300 477062 323534 477788
rect 322344 475098 323534 477062
rect 322344 474174 322604 475098
rect 323280 474174 323534 475098
rect 322344 473894 323534 474174
rect 412344 477788 413534 477990
rect 412344 477062 412608 477788
rect 413300 477062 413534 477788
rect 412344 475098 413534 477062
rect 412344 474174 412604 475098
rect 413280 474174 413534 475098
rect 412344 473894 413534 474174
rect 502344 477788 503534 477990
rect 502344 477062 502608 477788
rect 503300 477062 503534 477788
rect 502344 475098 503534 477062
rect 502344 474174 502604 475098
rect 503280 474174 503534 475098
rect 502344 473894 503534 474174
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 64524 389424 65714 389832
rect 64524 388500 64750 389424
rect 65426 388500 65714 389424
rect 64524 386810 65714 388500
rect 64524 386084 64790 386810
rect 65482 386084 65714 386810
rect 64524 385736 65714 386084
rect 154524 389424 155714 389832
rect 154524 388500 154750 389424
rect 155426 388500 155714 389424
rect 154524 386810 155714 388500
rect 154524 386084 154790 386810
rect 155482 386084 155714 386810
rect 154524 385736 155714 386084
rect 244524 389424 245714 389832
rect 244524 388500 244750 389424
rect 245426 388500 245714 389424
rect 244524 386810 245714 388500
rect 244524 386084 244790 386810
rect 245482 386084 245714 386810
rect 244524 385736 245714 386084
rect 334524 389424 335714 389832
rect 334524 388500 334750 389424
rect 335426 388500 335714 389424
rect 334524 386810 335714 388500
rect 334524 386084 334790 386810
rect 335482 386084 335714 386810
rect 334524 385736 335714 386084
rect 424524 389424 425714 389832
rect 424524 388500 424750 389424
rect 425426 388500 425714 389424
rect 424524 386810 425714 388500
rect 424524 386084 424790 386810
rect 425482 386084 425714 386810
rect 424524 385736 425714 386084
rect 514524 389424 515714 389832
rect 514524 388500 514750 389424
rect 515426 388500 515714 389424
rect 514524 386810 515714 388500
rect 514524 386084 514790 386810
rect 515482 386084 515714 386810
rect 514524 385736 515714 386084
rect -800 381864 480 381976
rect 57138 381380 58098 381620
rect -800 380682 480 380794
rect 57138 380600 57318 381380
rect 57978 380600 58098 381380
rect 57138 379935 58098 380600
rect -800 379500 480 379612
rect 57138 379190 57278 379935
rect 57958 379190 58098 379935
rect 57138 378735 58098 379190
rect 60858 381380 61818 381620
rect 60858 380600 61038 381380
rect 61698 380600 61818 381380
rect 60858 379965 61818 380600
rect 60858 379220 60998 379965
rect 61678 379220 61818 379965
rect 60858 378735 61818 379220
rect 147138 381380 148098 381620
rect 147138 380600 147318 381380
rect 147978 380600 148098 381380
rect 147138 379935 148098 380600
rect 147138 379190 147278 379935
rect 147958 379190 148098 379935
rect 147138 378735 148098 379190
rect 150858 381380 151818 381620
rect 150858 380600 151038 381380
rect 151698 380600 151818 381380
rect 150858 379965 151818 380600
rect 150858 379220 150998 379965
rect 151678 379220 151818 379965
rect 150858 378735 151818 379220
rect 237138 381380 238098 381620
rect 237138 380600 237318 381380
rect 237978 380600 238098 381380
rect -800 378318 480 378430
rect 237138 378380 238098 380600
rect 237138 377720 237318 378380
rect 237978 377720 238098 378380
rect 237138 377540 238098 377720
rect 240858 381380 241818 381620
rect 240858 380600 241038 381380
rect 241698 380600 241818 381380
rect 240858 378380 241818 380600
rect 240858 377720 241038 378380
rect 241698 377720 241818 378380
rect 240858 377540 241818 377720
rect 327138 381380 328098 381620
rect 327138 380600 327318 381380
rect 327978 380600 328098 381380
rect 327138 378380 328098 380600
rect 327138 377720 327318 378380
rect 327978 377720 328098 378380
rect 327138 377540 328098 377720
rect 330858 381380 331818 381620
rect 330858 380600 331038 381380
rect 331698 380600 331818 381380
rect 330858 378380 331818 380600
rect 330858 377720 331038 378380
rect 331698 377720 331818 378380
rect 330858 377540 331818 377720
rect 417138 381380 418098 381620
rect 417138 380600 417318 381380
rect 417978 380600 418098 381380
rect 417138 378380 418098 380600
rect 417138 377720 417318 378380
rect 417978 377720 418098 378380
rect 417138 377540 418098 377720
rect 420858 381380 421818 381620
rect 420858 380600 421038 381380
rect 421698 380600 421818 381380
rect 420858 378380 421818 380600
rect 420858 377720 421038 378380
rect 421698 377720 421818 378380
rect 420858 377540 421818 377720
rect 507138 381380 508098 381620
rect 507138 380600 507318 381380
rect 507978 380600 508098 381380
rect 507138 378380 508098 380600
rect 507138 377720 507318 378380
rect 507978 377720 508098 378380
rect 507138 377540 508098 377720
rect 510858 381380 511818 381620
rect 510858 380600 511038 381380
rect 511698 380600 511818 381380
rect 510858 378380 511818 380600
rect 510858 377720 511038 378380
rect 511698 377720 511818 378380
rect 510858 377540 511818 377720
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 230428 374443 231386 374448
rect 229045 373495 229051 374443
rect 229999 373495 230433 374443
rect 231381 373495 231386 374443
rect 230428 373490 231386 373495
rect 320958 372354 321294 372359
rect 320269 372028 320275 372354
rect 320601 372028 320963 372354
rect 321289 372028 321294 372354
rect 320958 372023 321294 372028
rect 339786 371700 340218 371705
rect 339786 371278 339791 371700
rect 340213 371278 340369 371700
rect 340791 371278 340797 371700
rect 415834 371300 417066 372058
rect 417542 371794 417798 371830
rect 423771 371821 424645 371841
rect 417542 371668 417598 371794
rect 417746 371668 417798 371794
rect 339786 371273 340218 371278
rect 415834 371100 415884 371300
rect 416084 371294 417284 371300
rect 417542 371294 417798 371668
rect 423278 371540 424645 371821
rect 423278 371486 423948 371540
rect 416084 371100 417798 371294
rect 422664 371408 423948 371486
rect 422664 371204 422700 371408
rect 422830 371204 423948 371408
rect 422664 371172 423948 371204
rect 415834 370750 417066 371100
rect 417216 371094 417798 371100
rect 417542 371092 417798 371094
rect 423278 371090 423948 371172
rect 424398 371090 424645 371540
rect 423278 370805 424645 371090
rect 505834 371300 507066 372058
rect 511638 371940 511858 371960
rect 511638 371780 511658 371940
rect 511818 371938 511858 371940
rect 511818 371821 512975 371938
rect 513771 371821 514645 371841
rect 511818 371784 514645 371821
rect 511818 371780 511858 371784
rect 511638 371760 511858 371780
rect 512821 371540 514645 371784
rect 505834 371100 505884 371300
rect 506084 371260 507798 371300
rect 506084 371140 507558 371260
rect 507758 371140 507798 371260
rect 512821 371255 513948 371540
rect 506084 371100 507798 371140
rect 505834 370750 507066 371100
rect 512817 371090 513948 371255
rect 514398 371090 514645 371540
rect 512817 370805 514645 371090
rect 49658 369730 50758 369735
rect 49658 368640 49663 369730
rect 50753 368640 50758 369730
rect 139658 369730 140758 369735
rect 49658 368635 50758 368640
rect 68313 369300 69193 369305
rect 49663 367805 50753 368635
rect 68313 368430 68318 369300
rect 69188 368430 69193 369300
rect 139658 368640 139663 369730
rect 140753 368640 140758 369730
rect 139658 368635 140758 368640
rect 158313 369300 159193 369305
rect 68313 368425 69193 368430
rect 49663 366709 50753 366715
rect 68318 367410 69188 368425
rect 139663 367805 140753 368635
rect 158313 368430 158318 369300
rect 159188 368430 159193 369300
rect 158313 368425 159193 368430
rect 139663 366709 140753 366715
rect 158318 367410 159188 368425
rect 68318 366534 69188 366540
rect 247586 368089 249097 368093
rect 247586 368088 249825 368089
rect 247586 366587 247591 368088
rect 249092 366588 249825 368088
rect 251326 366588 251332 368089
rect 249092 366587 249097 366588
rect 247586 366582 249097 366587
rect 158318 366534 159188 366540
rect 237078 365900 238038 366080
rect 57073 365130 58033 365275
rect 57073 364385 57193 365130
rect 57873 364665 58033 365130
rect 60798 365130 61758 365220
rect 57873 364385 58038 364665
rect 57073 364315 58038 364385
rect 57078 363020 58038 364315
rect 57078 362240 57258 363020
rect 57918 362240 58038 363020
rect 57078 362000 58038 362240
rect 60798 364385 60963 365130
rect 61643 364385 61758 365130
rect 60798 363020 61758 364385
rect 147073 365130 148033 365275
rect 237078 365240 237258 365900
rect 237918 365240 238038 365900
rect 147073 364385 147193 365130
rect 147873 364665 148033 365130
rect 150798 365130 151758 365220
rect 147873 364385 148038 364665
rect 147073 364315 148038 364385
rect 60798 362240 60978 363020
rect 61638 362240 61758 363020
rect 60798 362000 61758 362240
rect 147078 363020 148038 364315
rect 147078 362240 147258 363020
rect 147918 362240 148038 363020
rect 147078 362000 148038 362240
rect 150798 364385 150963 365130
rect 151643 364385 151758 365130
rect 150798 363020 151758 364385
rect 150798 362240 150978 363020
rect 151638 362240 151758 363020
rect 150798 362000 151758 362240
rect 237078 363020 238038 365240
rect 237078 362240 237258 363020
rect 237918 362240 238038 363020
rect 237078 362000 238038 362240
rect 240798 365900 241758 366080
rect 240798 365240 240978 365900
rect 241638 365240 241758 365900
rect 240798 363020 241758 365240
rect 240798 362240 240978 363020
rect 241638 362240 241758 363020
rect 240798 362000 241758 362240
rect 327078 365900 328038 366080
rect 327078 365240 327258 365900
rect 327918 365240 328038 365900
rect 327078 363020 328038 365240
rect 327078 362240 327258 363020
rect 327918 362240 328038 363020
rect 327078 362000 328038 362240
rect 330798 365900 331758 366080
rect 330798 365240 330978 365900
rect 331638 365240 331758 365900
rect 330798 363020 331758 365240
rect 330798 362240 330978 363020
rect 331638 362240 331758 363020
rect 330798 362000 331758 362240
rect 417078 365900 418038 366080
rect 417078 365240 417258 365900
rect 417918 365240 418038 365900
rect 417078 363020 418038 365240
rect 417078 362240 417258 363020
rect 417918 362240 418038 363020
rect 417078 362000 418038 362240
rect 420798 365900 421758 366080
rect 420798 365240 420978 365900
rect 421638 365240 421758 365900
rect 420798 363020 421758 365240
rect 420798 362240 420978 363020
rect 421638 362240 421758 363020
rect 420798 362000 421758 362240
rect 507078 365900 508038 366080
rect 507078 365240 507258 365900
rect 507918 365240 508038 365900
rect 507078 363020 508038 365240
rect 507078 362240 507258 363020
rect 507918 362240 508038 363020
rect 507078 362000 508038 362240
rect 510798 365900 511758 366080
rect 510798 365240 510978 365900
rect 511638 365240 511758 365900
rect 510798 363020 511758 365240
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 510798 362240 510978 363020
rect 511638 362240 511758 363020
rect 583520 362420 584800 362532
rect 510798 362000 511758 362240
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect 52344 357788 53534 357990
rect 52344 357062 52608 357788
rect 53300 357062 53534 357788
rect 52344 355098 53534 357062
rect 52344 354174 52604 355098
rect 53280 354174 53534 355098
rect 52344 353894 53534 354174
rect 142344 357788 143534 357990
rect 142344 357062 142608 357788
rect 143300 357062 143534 357788
rect 142344 355098 143534 357062
rect 142344 354174 142604 355098
rect 143280 354174 143534 355098
rect 142344 353894 143534 354174
rect 232344 357788 233534 357990
rect 232344 357062 232608 357788
rect 233300 357062 233534 357788
rect 232344 355098 233534 357062
rect 232344 354174 232604 355098
rect 233280 354174 233534 355098
rect 232344 353894 233534 354174
rect 322344 357788 323534 357990
rect 322344 357062 322608 357788
rect 323300 357062 323534 357788
rect 322344 355098 323534 357062
rect 322344 354174 322604 355098
rect 323280 354174 323534 355098
rect 322344 353894 323534 354174
rect 412344 357788 413534 357990
rect 412344 357062 412608 357788
rect 413300 357062 413534 357788
rect 412344 355098 413534 357062
rect 412344 354174 412604 355098
rect 413280 354174 413534 355098
rect 412344 353894 413534 354174
rect 502344 357788 503534 357990
rect 502344 357062 502608 357788
rect 503300 357062 503534 357788
rect 502344 355098 503534 357062
rect 502344 354174 502604 355098
rect 503280 354174 503534 355098
rect 502344 353894 503534 354174
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 64524 269424 65714 269832
rect 64524 268500 64750 269424
rect 65426 268500 65714 269424
rect 64524 266810 65714 268500
rect 64524 266084 64790 266810
rect 65482 266084 65714 266810
rect 64524 265736 65714 266084
rect 153648 269220 154838 269628
rect 153648 268296 153874 269220
rect 154550 268296 154838 269220
rect 153648 266606 154838 268296
rect 153648 265880 153914 266606
rect 154606 265880 154838 266606
rect 153648 265532 154838 265880
rect 244902 269032 246092 269440
rect 244902 268108 245128 269032
rect 245804 268108 246092 269032
rect 244902 266418 246092 268108
rect 244902 265692 245168 266418
rect 245860 265692 246092 266418
rect 334524 269424 335714 269832
rect 334524 268500 334750 269424
rect 335426 268500 335714 269424
rect 334524 266810 335714 268500
rect 334524 266084 334790 266810
rect 335482 266084 335714 266810
rect 334524 265736 335714 266084
rect 424524 269424 425714 269832
rect 424524 268500 424750 269424
rect 425426 268500 425714 269424
rect 424524 266810 425714 268500
rect 424524 266084 424790 266810
rect 425482 266084 425714 266810
rect 424524 265736 425714 266084
rect 514524 269424 515714 269832
rect 514524 268500 514750 269424
rect 515426 268500 515714 269424
rect 583520 269230 584800 269342
rect 514524 266810 515714 268500
rect 514524 266084 514790 266810
rect 515482 266084 515714 266810
rect 514524 265736 515714 266084
rect 244902 265344 246092 265692
rect 57138 261380 58098 261620
rect 57138 260600 57318 261380
rect 57978 260600 58098 261380
rect 57138 258380 58098 260600
rect 57138 257720 57318 258380
rect 57978 257720 58098 258380
rect 57138 257540 58098 257720
rect 60858 261380 61818 261620
rect 60858 260600 61038 261380
rect 61698 260600 61818 261380
rect 60858 258380 61818 260600
rect 60858 257720 61038 258380
rect 61698 257720 61818 258380
rect 60858 257540 61818 257720
rect 146262 261176 147222 261416
rect 146262 260396 146442 261176
rect 147102 260396 147222 261176
rect 146262 258176 147222 260396
rect 146262 257516 146442 258176
rect 147102 257516 147222 258176
rect 146262 257336 147222 257516
rect 149982 261176 150942 261416
rect 327138 261380 328098 261620
rect 149982 260396 150162 261176
rect 150822 260396 150942 261176
rect 149982 258176 150942 260396
rect 149982 257516 150162 258176
rect 150822 257516 150942 258176
rect 149982 257336 150942 257516
rect 237516 260988 238476 261228
rect 237516 260208 237696 260988
rect 238356 260208 238476 260988
rect 237516 257988 238476 260208
rect 237516 257328 237696 257988
rect 238356 257328 238476 257988
rect 237516 257148 238476 257328
rect 241236 260988 242196 261228
rect 241236 260208 241416 260988
rect 242076 260208 242196 260988
rect 241236 257988 242196 260208
rect 241236 257328 241416 257988
rect 242076 257328 242196 257988
rect 327138 260600 327318 261380
rect 327978 260600 328098 261380
rect 327138 258380 328098 260600
rect 327138 257720 327318 258380
rect 327978 257720 328098 258380
rect 327138 257540 328098 257720
rect 330858 261380 331818 261620
rect 330858 260600 331038 261380
rect 331698 260600 331818 261380
rect 330858 258380 331818 260600
rect 417138 261380 418098 261620
rect 417138 260600 417318 261380
rect 417978 260600 418098 261380
rect 417138 259935 418098 260600
rect 417138 259190 417278 259935
rect 417958 259190 418098 259935
rect 417138 258735 418098 259190
rect 420858 261380 421818 261620
rect 420858 260600 421038 261380
rect 421698 260600 421818 261380
rect 420858 259965 421818 260600
rect 420858 259220 420998 259965
rect 421678 259220 421818 259965
rect 420858 258735 421818 259220
rect 507138 261380 508098 261620
rect 507138 260600 507318 261380
rect 507978 260600 508098 261380
rect 507138 259935 508098 260600
rect 507138 259190 507278 259935
rect 507958 259190 508098 259935
rect 507138 258735 508098 259190
rect 510858 261380 511818 261620
rect 510858 260600 511038 261380
rect 511698 260600 511818 261380
rect 510858 259965 511818 260600
rect 510858 259220 510998 259965
rect 511678 259220 511818 259965
rect 510858 258735 511818 259220
rect 330858 257720 331038 258380
rect 331698 257720 331818 258380
rect 330858 257540 331818 257720
rect 241236 257148 242196 257328
rect 320428 254443 321386 254448
rect 319045 253495 319051 254443
rect 319999 253495 320433 254443
rect 321381 253495 321386 254443
rect 320428 253490 321386 253495
rect -800 252398 480 252510
rect -800 251216 480 251328
rect 55834 251300 57066 252058
rect 231336 251962 231672 251967
rect 61638 251940 61858 251960
rect 61638 251780 61658 251940
rect 61818 251938 61858 251940
rect 61818 251821 62975 251938
rect 63771 251821 64645 251841
rect 61818 251784 64645 251821
rect 61818 251780 61858 251784
rect 61638 251760 61858 251780
rect 62821 251540 64645 251784
rect 55834 251100 55884 251300
rect 56084 251260 57798 251300
rect 56084 251140 57558 251260
rect 57758 251140 57798 251260
rect 62821 251255 63948 251540
rect 56084 251100 57798 251140
rect 55834 250750 57066 251100
rect 62817 251090 63948 251255
rect 64398 251090 64645 251540
rect 62817 250805 64645 251090
rect 144958 251096 146190 251854
rect 146666 251590 146922 251626
rect 152895 251617 153769 251637
rect 230647 251636 230653 251962
rect 230979 251636 231341 251962
rect 231667 251636 231672 251962
rect 231336 251631 231672 251636
rect 146666 251464 146722 251590
rect 146870 251464 146922 251590
rect 144958 250896 145008 251096
rect 145208 251090 146408 251096
rect 146666 251090 146922 251464
rect 152402 251336 153769 251617
rect 152402 251282 153072 251336
rect 145208 250896 146922 251090
rect 151788 251204 153072 251282
rect 151788 251000 151824 251204
rect 151954 251000 153072 251204
rect 151788 250968 153072 251000
rect 144958 250546 146190 250896
rect 146340 250890 146922 250896
rect 146666 250888 146922 250890
rect 152402 250886 153072 250968
rect 153522 250886 153769 251336
rect 152402 250601 153769 250886
rect 250164 251308 250596 251313
rect 250164 250886 250169 251308
rect 250591 250886 250747 251308
rect 251169 250886 251175 251308
rect 250164 250881 250596 250886
rect -800 250034 480 250146
rect 409658 249730 410758 249735
rect -800 248852 480 248964
rect 409658 248640 409663 249730
rect 410753 248640 410758 249730
rect 499658 249730 500758 249735
rect 409658 248635 410758 248640
rect 428313 249300 429193 249305
rect 337586 248089 339097 248093
rect 337586 248088 339825 248089
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 337586 246587 337591 248088
rect 339092 246588 339825 248088
rect 341326 246588 341332 248089
rect 409663 247805 410753 248635
rect 428313 248430 428318 249300
rect 429188 248430 429193 249300
rect 499658 248640 499663 249730
rect 500753 248640 500758 249730
rect 499658 248635 500758 248640
rect 518313 249300 519193 249305
rect 428313 248425 429193 248430
rect 409663 246709 410753 246715
rect 428318 247410 429188 248425
rect 339092 246587 339097 246588
rect 337586 246582 339097 246587
rect 499663 247805 500753 248635
rect 518313 248430 518318 249300
rect 519188 248430 519193 249300
rect 518313 248425 519193 248430
rect 499663 246709 500753 246715
rect 518318 247410 519188 248425
rect 428318 246534 429188 246540
rect 518318 246534 519188 246540
rect 57078 245900 58038 246080
rect 57078 245240 57258 245900
rect 57918 245240 58038 245900
rect 57078 243020 58038 245240
rect 57078 242240 57258 243020
rect 57918 242240 58038 243020
rect 57078 242000 58038 242240
rect 60798 245900 61758 246080
rect 60798 245240 60978 245900
rect 61638 245240 61758 245900
rect 327078 245900 328038 246080
rect 60798 243020 61758 245240
rect 60798 242240 60978 243020
rect 61638 242240 61758 243020
rect 60798 242000 61758 242240
rect 146202 245696 147162 245876
rect 146202 245036 146382 245696
rect 147042 245036 147162 245696
rect 146202 242816 147162 245036
rect 146202 242036 146382 242816
rect 147042 242036 147162 242816
rect 146202 241796 147162 242036
rect 149922 245696 150882 245876
rect 149922 245036 150102 245696
rect 150762 245036 150882 245696
rect 149922 242816 150882 245036
rect 149922 242036 150102 242816
rect 150762 242036 150882 242816
rect 149922 241796 150882 242036
rect 237456 245508 238416 245688
rect 237456 244848 237636 245508
rect 238296 244848 238416 245508
rect 237456 242628 238416 244848
rect 237456 241848 237636 242628
rect 238296 241848 238416 242628
rect 237456 241608 238416 241848
rect 241176 245508 242136 245688
rect 241176 244848 241356 245508
rect 242016 244848 242136 245508
rect 241176 242628 242136 244848
rect 241176 241848 241356 242628
rect 242016 241848 242136 242628
rect 327078 245240 327258 245900
rect 327918 245240 328038 245900
rect 327078 243020 328038 245240
rect 327078 242240 327258 243020
rect 327918 242240 328038 243020
rect 327078 242000 328038 242240
rect 330798 245900 331758 246080
rect 330798 245240 330978 245900
rect 331638 245240 331758 245900
rect 330798 243020 331758 245240
rect 417073 245130 418033 245275
rect 417073 244385 417193 245130
rect 417873 244665 418033 245130
rect 420798 245130 421758 245220
rect 417873 244385 418038 244665
rect 417073 244315 418038 244385
rect 330798 242240 330978 243020
rect 331638 242240 331758 243020
rect 330798 242000 331758 242240
rect 417078 243020 418038 244315
rect 417078 242240 417258 243020
rect 417918 242240 418038 243020
rect 417078 242000 418038 242240
rect 420798 244385 420963 245130
rect 421643 244385 421758 245130
rect 420798 243020 421758 244385
rect 507073 245130 508033 245275
rect 507073 244385 507193 245130
rect 507873 244665 508033 245130
rect 510798 245130 511758 245220
rect 507873 244385 508038 244665
rect 507073 244315 508038 244385
rect 420798 242240 420978 243020
rect 421638 242240 421758 243020
rect 420798 242000 421758 242240
rect 507078 243020 508038 244315
rect 507078 242240 507258 243020
rect 507918 242240 508038 243020
rect 507078 242000 508038 242240
rect 510798 244385 510963 245130
rect 511643 244385 511758 245130
rect 510798 243020 511758 244385
rect 510798 242240 510978 243020
rect 511638 242240 511758 243020
rect 510798 242000 511758 242240
rect 241176 241608 242136 241848
rect 52344 237788 53534 237990
rect 52344 237062 52608 237788
rect 53300 237062 53534 237788
rect 322344 237788 323534 237990
rect 52344 235098 53534 237062
rect 52344 234174 52604 235098
rect 53280 234174 53534 235098
rect 52344 233894 53534 234174
rect 141468 237584 142658 237786
rect 141468 236858 141732 237584
rect 142424 236858 142658 237584
rect 141468 234894 142658 236858
rect 141468 233970 141728 234894
rect 142404 233970 142658 234894
rect 141468 233690 142658 233970
rect 232722 237396 233912 237598
rect 232722 236670 232986 237396
rect 233678 236670 233912 237396
rect 232722 234706 233912 236670
rect 232722 233782 232982 234706
rect 233658 233782 233912 234706
rect 322344 237062 322608 237788
rect 323300 237062 323534 237788
rect 322344 235098 323534 237062
rect 322344 234174 322604 235098
rect 323280 234174 323534 235098
rect 322344 233894 323534 234174
rect 412344 237788 413534 237990
rect 412344 237062 412608 237788
rect 413300 237062 413534 237788
rect 412344 235098 413534 237062
rect 412344 234174 412604 235098
rect 413280 234174 413534 235098
rect 412344 233894 413534 234174
rect 502344 237788 503534 237990
rect 502344 237062 502608 237788
rect 503300 237062 503534 237788
rect 502344 235098 503534 237062
rect 582340 235230 584800 240030
rect 502344 234174 502604 235098
rect 503280 234174 503534 235098
rect 502344 233894 503534 234174
rect 232722 233502 233912 233782
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 57138 155280 58098 155520
rect 57138 154500 57318 155280
rect 57978 154500 58098 155280
rect 57138 152280 58098 154500
rect 57138 151620 57318 152280
rect 57978 151620 58098 152280
rect 57138 151440 58098 151620
rect 60858 155280 61818 155520
rect 60858 154500 61038 155280
rect 61698 154500 61818 155280
rect 60858 152280 61818 154500
rect 60858 151620 61038 152280
rect 61698 151620 61818 152280
rect 60858 151440 61818 151620
rect 147138 155280 148098 155520
rect 147138 154500 147318 155280
rect 147978 154500 148098 155280
rect 147138 152280 148098 154500
rect 147138 151620 147318 152280
rect 147978 151620 148098 152280
rect 147138 151440 148098 151620
rect 150858 155280 151818 155520
rect 150858 154500 151038 155280
rect 151698 154500 151818 155280
rect 150858 152280 151818 154500
rect 150858 151620 151038 152280
rect 151698 151620 151818 152280
rect 150858 151440 151818 151620
rect 237138 155280 238098 155520
rect 237138 154500 237318 155280
rect 237978 154500 238098 155280
rect 237138 152280 238098 154500
rect 237138 151620 237318 152280
rect 237978 151620 238098 152280
rect 237138 151440 238098 151620
rect 240858 155280 241818 155520
rect 240858 154500 241038 155280
rect 241698 154500 241818 155280
rect 240858 152280 241818 154500
rect 240858 151620 241038 152280
rect 241698 151620 241818 152280
rect 240858 151440 241818 151620
rect 327138 155280 328098 155520
rect 327138 154500 327318 155280
rect 327978 154500 328098 155280
rect 327138 152280 328098 154500
rect 327138 151620 327318 152280
rect 327978 151620 328098 152280
rect 327138 151440 328098 151620
rect 330858 155280 331818 155520
rect 330858 154500 331038 155280
rect 331698 154500 331818 155280
rect 330858 152280 331818 154500
rect 330858 151620 331038 152280
rect 331698 151620 331818 152280
rect 330858 151440 331818 151620
rect 417138 155280 418098 155520
rect 417138 154500 417318 155280
rect 417978 154500 418098 155280
rect 417138 152280 418098 154500
rect 417138 151620 417318 152280
rect 417978 151620 418098 152280
rect 417138 151440 418098 151620
rect 420858 155280 421818 155520
rect 420858 154500 421038 155280
rect 421698 154500 421818 155280
rect 420858 152280 421818 154500
rect 420858 151620 421038 152280
rect 421698 151620 421818 152280
rect 420858 151440 421818 151620
rect 507138 155280 508098 155520
rect 507138 154500 507318 155280
rect 507978 154500 508098 155280
rect 507138 152280 508098 154500
rect 507138 151620 507318 152280
rect 507978 151620 508098 152280
rect 507138 151440 508098 151620
rect 510858 155280 511818 155520
rect 510858 154500 511038 155280
rect 511698 154500 511818 155280
rect 510858 152280 511818 154500
rect 510858 151620 511038 152280
rect 511698 151620 511818 152280
rect 510858 151440 511818 151620
rect 582340 146830 584800 151630
rect 55834 145200 57066 145958
rect 61638 145840 61858 145860
rect 61638 145680 61658 145840
rect 61818 145838 61858 145840
rect 61818 145721 62975 145838
rect 63771 145721 64645 145741
rect 61818 145684 64645 145721
rect 61818 145680 61858 145684
rect 61638 145660 61858 145680
rect 62821 145440 64645 145684
rect 55834 145000 55884 145200
rect 56084 145160 57798 145200
rect 56084 145040 57558 145160
rect 57758 145040 57798 145160
rect 62821 145155 63948 145440
rect 56084 145000 57798 145040
rect 55834 144650 57066 145000
rect 62817 144990 63948 145155
rect 64398 144990 64645 145440
rect 62817 144705 64645 144990
rect 145834 145200 147066 145958
rect 151638 145840 151858 145860
rect 151638 145680 151658 145840
rect 151818 145838 151858 145840
rect 151818 145721 152975 145838
rect 153771 145721 154645 145741
rect 151818 145684 154645 145721
rect 151818 145680 151858 145684
rect 151638 145660 151858 145680
rect 152821 145440 154645 145684
rect 145834 145000 145884 145200
rect 146084 145160 147798 145200
rect 146084 145040 147558 145160
rect 147758 145040 147798 145160
rect 152821 145155 153948 145440
rect 146084 145000 147798 145040
rect 145834 144650 147066 145000
rect 152817 144990 153948 145155
rect 154398 144990 154645 145440
rect 152817 144705 154645 144990
rect 235834 145200 237066 145958
rect 241638 145840 241858 145860
rect 241638 145680 241658 145840
rect 241818 145838 241858 145840
rect 241818 145721 242975 145838
rect 243771 145721 244645 145741
rect 241818 145684 244645 145721
rect 241818 145680 241858 145684
rect 241638 145660 241858 145680
rect 242821 145440 244645 145684
rect 235834 145000 235884 145200
rect 236084 145160 237798 145200
rect 236084 145040 237558 145160
rect 237758 145040 237798 145160
rect 242821 145155 243948 145440
rect 236084 145000 237798 145040
rect 235834 144650 237066 145000
rect 242817 144990 243948 145155
rect 244398 144990 244645 145440
rect 242817 144705 244645 144990
rect 325834 145200 327066 145958
rect 331638 145840 331858 145860
rect 331638 145680 331658 145840
rect 331818 145838 331858 145840
rect 331818 145721 332975 145838
rect 333771 145721 334645 145741
rect 331818 145684 334645 145721
rect 331818 145680 331858 145684
rect 331638 145660 331858 145680
rect 332821 145440 334645 145684
rect 325834 145000 325884 145200
rect 326084 145160 327798 145200
rect 326084 145040 327558 145160
rect 327758 145040 327798 145160
rect 332821 145155 333948 145440
rect 326084 145000 327798 145040
rect 325834 144650 327066 145000
rect 332817 144990 333948 145155
rect 334398 144990 334645 145440
rect 332817 144705 334645 144990
rect 415834 145200 417066 145958
rect 421638 145840 421858 145860
rect 421638 145680 421658 145840
rect 421818 145838 421858 145840
rect 421818 145721 422975 145838
rect 423771 145721 424645 145741
rect 421818 145684 424645 145721
rect 421818 145680 421858 145684
rect 421638 145660 421858 145680
rect 422821 145440 424645 145684
rect 415834 145000 415884 145200
rect 416084 145160 417798 145200
rect 416084 145040 417558 145160
rect 417758 145040 417798 145160
rect 422821 145155 423948 145440
rect 416084 145000 417798 145040
rect 415834 144650 417066 145000
rect 422817 144990 423948 145155
rect 424398 144990 424645 145440
rect 422817 144705 424645 144990
rect 505834 145200 507066 145958
rect 511638 145840 511858 145860
rect 511638 145680 511658 145840
rect 511818 145838 511858 145840
rect 511818 145721 512975 145838
rect 513771 145721 514645 145741
rect 511818 145684 514645 145721
rect 511818 145680 511858 145684
rect 511638 145660 511858 145680
rect 512821 145440 514645 145684
rect 505834 145000 505884 145200
rect 506084 145160 507798 145200
rect 506084 145040 507558 145160
rect 507758 145040 507798 145160
rect 512821 145155 513948 145440
rect 506084 145000 507798 145040
rect 505834 144650 507066 145000
rect 512817 144990 513948 145155
rect 514398 144990 514645 145440
rect 512817 144705 514645 144990
rect 57078 139800 58038 139980
rect 57078 139140 57258 139800
rect 57918 139140 58038 139800
rect 57078 136920 58038 139140
rect 57078 136140 57258 136920
rect 57918 136140 58038 136920
rect 57078 135900 58038 136140
rect 60798 139800 61758 139980
rect 60798 139140 60978 139800
rect 61638 139140 61758 139800
rect 60798 136920 61758 139140
rect 60798 136140 60978 136920
rect 61638 136140 61758 136920
rect 60798 135900 61758 136140
rect 147078 139800 148038 139980
rect 147078 139140 147258 139800
rect 147918 139140 148038 139800
rect 147078 136920 148038 139140
rect 147078 136140 147258 136920
rect 147918 136140 148038 136920
rect 147078 135900 148038 136140
rect 150798 139800 151758 139980
rect 150798 139140 150978 139800
rect 151638 139140 151758 139800
rect 150798 136920 151758 139140
rect 150798 136140 150978 136920
rect 151638 136140 151758 136920
rect 150798 135900 151758 136140
rect 237078 139800 238038 139980
rect 237078 139140 237258 139800
rect 237918 139140 238038 139800
rect 237078 136920 238038 139140
rect 237078 136140 237258 136920
rect 237918 136140 238038 136920
rect 237078 135900 238038 136140
rect 240798 139800 241758 139980
rect 240798 139140 240978 139800
rect 241638 139140 241758 139800
rect 240798 136920 241758 139140
rect 240798 136140 240978 136920
rect 241638 136140 241758 136920
rect 240798 135900 241758 136140
rect 327078 139800 328038 139980
rect 327078 139140 327258 139800
rect 327918 139140 328038 139800
rect 327078 136920 328038 139140
rect 327078 136140 327258 136920
rect 327918 136140 328038 136920
rect 327078 135900 328038 136140
rect 330798 139800 331758 139980
rect 330798 139140 330978 139800
rect 331638 139140 331758 139800
rect 330798 136920 331758 139140
rect 330798 136140 330978 136920
rect 331638 136140 331758 136920
rect 330798 135900 331758 136140
rect 417078 139800 418038 139980
rect 417078 139140 417258 139800
rect 417918 139140 418038 139800
rect 417078 136920 418038 139140
rect 417078 136140 417258 136920
rect 417918 136140 418038 136920
rect 417078 135900 418038 136140
rect 420798 139800 421758 139980
rect 420798 139140 420978 139800
rect 421638 139140 421758 139800
rect 420798 136920 421758 139140
rect 420798 136140 420978 136920
rect 421638 136140 421758 136920
rect 420798 135900 421758 136140
rect 507078 139800 508038 139980
rect 507078 139140 507258 139800
rect 507918 139140 508038 139800
rect 507078 136920 508038 139140
rect 507078 136140 507258 136920
rect 507918 136140 508038 136920
rect 507078 135900 508038 136140
rect 510798 139800 511758 139980
rect 510798 139140 510978 139800
rect 511638 139140 511758 139800
rect 510798 136920 511758 139140
rect 510798 136140 510978 136920
rect 511638 136140 511758 136920
rect 582340 136830 584800 141630
rect 510798 135900 511758 136140
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 57138 65280 58098 65520
rect 57138 64500 57318 65280
rect 57978 64500 58098 65280
rect 57138 62280 58098 64500
rect 57138 61620 57318 62280
rect 57978 61620 58098 62280
rect 57138 61440 58098 61620
rect 60858 65280 61818 65520
rect 60858 64500 61038 65280
rect 61698 64500 61818 65280
rect 60858 62280 61818 64500
rect 60858 61620 61038 62280
rect 61698 61620 61818 62280
rect 60858 61440 61818 61620
rect 147138 65280 148098 65520
rect 147138 64500 147318 65280
rect 147978 64500 148098 65280
rect 147138 62280 148098 64500
rect 147138 61620 147318 62280
rect 147978 61620 148098 62280
rect 147138 61440 148098 61620
rect 150858 65280 151818 65520
rect 150858 64500 151038 65280
rect 151698 64500 151818 65280
rect 150858 62280 151818 64500
rect 150858 61620 151038 62280
rect 151698 61620 151818 62280
rect 150858 61440 151818 61620
rect 237138 65280 238098 65520
rect 237138 64500 237318 65280
rect 237978 64500 238098 65280
rect 237138 62280 238098 64500
rect 237138 61620 237318 62280
rect 237978 61620 238098 62280
rect 237138 61440 238098 61620
rect 240858 65280 241818 65520
rect 240858 64500 241038 65280
rect 241698 64500 241818 65280
rect 240858 62280 241818 64500
rect 240858 61620 241038 62280
rect 241698 61620 241818 62280
rect 240858 61440 241818 61620
rect 327138 65280 328098 65520
rect 327138 64500 327318 65280
rect 327978 64500 328098 65280
rect 327138 62280 328098 64500
rect 327138 61620 327318 62280
rect 327978 61620 328098 62280
rect 327138 61440 328098 61620
rect 330858 65280 331818 65520
rect 330858 64500 331038 65280
rect 331698 64500 331818 65280
rect 330858 62280 331818 64500
rect 330858 61620 331038 62280
rect 331698 61620 331818 62280
rect 330858 61440 331818 61620
rect 417138 65280 418098 65520
rect 417138 64500 417318 65280
rect 417978 64500 418098 65280
rect 417138 62280 418098 64500
rect 417138 61620 417318 62280
rect 417978 61620 418098 62280
rect 417138 61440 418098 61620
rect 420858 65280 421818 65520
rect 420858 64500 421038 65280
rect 421698 64500 421818 65280
rect 420858 62280 421818 64500
rect 420858 61620 421038 62280
rect 421698 61620 421818 62280
rect 420858 61440 421818 61620
rect 507138 65280 508098 65520
rect 507138 64500 507318 65280
rect 507978 64500 508098 65280
rect 507138 62280 508098 64500
rect 507138 61620 507318 62280
rect 507978 61620 508098 62280
rect 507138 61440 508098 61620
rect 510858 65280 511818 65520
rect 510858 64500 511038 65280
rect 511698 64500 511818 65280
rect 510858 62280 511818 64500
rect 510858 61620 511038 62280
rect 511698 61620 511818 62280
rect 510858 61440 511818 61620
rect 55834 55200 57066 55958
rect 61638 55840 61858 55860
rect 61638 55680 61658 55840
rect 61818 55838 61858 55840
rect 61818 55721 62975 55838
rect 63771 55721 64645 55741
rect 61818 55684 64645 55721
rect 61818 55680 61858 55684
rect 61638 55660 61858 55680
rect 62821 55440 64645 55684
rect 55834 55000 55884 55200
rect 56084 55160 57798 55200
rect 56084 55040 57558 55160
rect 57758 55040 57798 55160
rect 62821 55155 63948 55440
rect 56084 55000 57798 55040
rect 55834 54650 57066 55000
rect 62817 54990 63948 55155
rect 64398 54990 64645 55440
rect 62817 54705 64645 54990
rect 145834 55200 147066 55958
rect 151638 55840 151858 55860
rect 151638 55680 151658 55840
rect 151818 55838 151858 55840
rect 151818 55721 152975 55838
rect 153771 55721 154645 55741
rect 151818 55684 154645 55721
rect 151818 55680 151858 55684
rect 151638 55660 151858 55680
rect 152821 55440 154645 55684
rect 145834 55000 145884 55200
rect 146084 55160 147798 55200
rect 146084 55040 147558 55160
rect 147758 55040 147798 55160
rect 152821 55155 153948 55440
rect 146084 55000 147798 55040
rect 145834 54650 147066 55000
rect 152817 54990 153948 55155
rect 154398 54990 154645 55440
rect 152817 54705 154645 54990
rect 235834 55200 237066 55958
rect 241638 55840 241858 55860
rect 241638 55680 241658 55840
rect 241818 55838 241858 55840
rect 241818 55721 242975 55838
rect 243771 55721 244645 55741
rect 241818 55684 244645 55721
rect 241818 55680 241858 55684
rect 241638 55660 241858 55680
rect 242821 55440 244645 55684
rect 235834 55000 235884 55200
rect 236084 55160 237798 55200
rect 236084 55040 237558 55160
rect 237758 55040 237798 55160
rect 242821 55155 243948 55440
rect 236084 55000 237798 55040
rect 235834 54650 237066 55000
rect 242817 54990 243948 55155
rect 244398 54990 244645 55440
rect 242817 54705 244645 54990
rect 325834 55200 327066 55958
rect 331638 55840 331858 55860
rect 331638 55680 331658 55840
rect 331818 55838 331858 55840
rect 331818 55721 332975 55838
rect 333771 55721 334645 55741
rect 331818 55684 334645 55721
rect 331818 55680 331858 55684
rect 331638 55660 331858 55680
rect 332821 55440 334645 55684
rect 325834 55000 325884 55200
rect 326084 55160 327798 55200
rect 326084 55040 327558 55160
rect 327758 55040 327798 55160
rect 332821 55155 333948 55440
rect 326084 55000 327798 55040
rect 325834 54650 327066 55000
rect 332817 54990 333948 55155
rect 334398 54990 334645 55440
rect 332817 54705 334645 54990
rect 415834 55200 417066 55958
rect 421638 55840 421858 55860
rect 421638 55680 421658 55840
rect 421818 55838 421858 55840
rect 421818 55721 422975 55838
rect 423771 55721 424645 55741
rect 421818 55684 424645 55721
rect 421818 55680 421858 55684
rect 421638 55660 421858 55680
rect 422821 55440 424645 55684
rect 415834 55000 415884 55200
rect 416084 55160 417798 55200
rect 416084 55040 417558 55160
rect 417758 55040 417798 55160
rect 422821 55155 423948 55440
rect 416084 55000 417798 55040
rect 415834 54650 417066 55000
rect 422817 54990 423948 55155
rect 424398 54990 424645 55440
rect 422817 54705 424645 54990
rect 505834 55200 507066 55958
rect 511638 55840 511858 55860
rect 511638 55680 511658 55840
rect 511818 55838 511858 55840
rect 511818 55721 512975 55838
rect 513771 55721 514645 55741
rect 511818 55684 514645 55721
rect 511818 55680 511858 55684
rect 511638 55660 511858 55680
rect 512821 55440 514645 55684
rect 505834 55000 505884 55200
rect 506084 55160 507798 55200
rect 506084 55040 507558 55160
rect 507758 55040 507798 55160
rect 512821 55155 513948 55440
rect 506084 55000 507798 55040
rect 505834 54650 507066 55000
rect 512817 54990 513948 55155
rect 514398 54990 514645 55440
rect 512817 54705 514645 54990
rect 583520 50460 584800 50572
rect 57078 49800 58038 49980
rect 57078 49140 57258 49800
rect 57918 49140 58038 49800
rect 57078 46920 58038 49140
rect 57078 46140 57258 46920
rect 57918 46140 58038 46920
rect 57078 45900 58038 46140
rect 60798 49800 61758 49980
rect 60798 49140 60978 49800
rect 61638 49140 61758 49800
rect 60798 46920 61758 49140
rect 60798 46140 60978 46920
rect 61638 46140 61758 46920
rect 60798 45900 61758 46140
rect 147078 49800 148038 49980
rect 147078 49140 147258 49800
rect 147918 49140 148038 49800
rect 147078 46920 148038 49140
rect 147078 46140 147258 46920
rect 147918 46140 148038 46920
rect 147078 45900 148038 46140
rect 150798 49800 151758 49980
rect 150798 49140 150978 49800
rect 151638 49140 151758 49800
rect 150798 46920 151758 49140
rect 150798 46140 150978 46920
rect 151638 46140 151758 46920
rect 150798 45900 151758 46140
rect 237078 49800 238038 49980
rect 237078 49140 237258 49800
rect 237918 49140 238038 49800
rect 237078 46920 238038 49140
rect 237078 46140 237258 46920
rect 237918 46140 238038 46920
rect 237078 45900 238038 46140
rect 240798 49800 241758 49980
rect 240798 49140 240978 49800
rect 241638 49140 241758 49800
rect 240798 46920 241758 49140
rect 240798 46140 240978 46920
rect 241638 46140 241758 46920
rect 240798 45900 241758 46140
rect 327078 49800 328038 49980
rect 327078 49140 327258 49800
rect 327918 49140 328038 49800
rect 327078 46920 328038 49140
rect 327078 46140 327258 46920
rect 327918 46140 328038 46920
rect 327078 45900 328038 46140
rect 330798 49800 331758 49980
rect 330798 49140 330978 49800
rect 331638 49140 331758 49800
rect 330798 46920 331758 49140
rect 330798 46140 330978 46920
rect 331638 46140 331758 46920
rect 330798 45900 331758 46140
rect 417078 49800 418038 49980
rect 417078 49140 417258 49800
rect 417918 49140 418038 49800
rect 417078 46920 418038 49140
rect 417078 46140 417258 46920
rect 417918 46140 418038 46920
rect 417078 45900 418038 46140
rect 420798 49800 421758 49980
rect 420798 49140 420978 49800
rect 421638 49140 421758 49800
rect 420798 46920 421758 49140
rect 420798 46140 420978 46920
rect 421638 46140 421758 46920
rect 420798 45900 421758 46140
rect 507078 49800 508038 49980
rect 507078 49140 507258 49800
rect 507918 49140 508038 49800
rect 507078 46920 508038 49140
rect 507078 46140 507258 46920
rect 507918 46140 508038 46920
rect 507078 45900 508038 46140
rect 510798 49800 511758 49980
rect 510798 49140 510978 49800
rect 511638 49140 511758 49800
rect 583520 49278 584800 49390
rect 510798 46920 511758 49140
rect 583520 48096 584800 48208
rect 510798 46140 510978 46920
rect 511638 46140 511758 46920
rect 583520 46914 584800 47026
rect 510798 45900 511758 46140
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 327120 666424 327780 667204
rect 57318 664500 57978 665280
rect 61038 664500 61698 665280
rect 147318 664500 147978 665280
rect 151038 664500 151698 665280
rect 237318 664500 237978 665280
rect 241038 664500 241698 665280
rect 330840 666424 331500 667204
rect 417120 666424 417780 667204
rect 420840 666424 421500 667204
rect 507120 666424 507780 667204
rect 510840 666424 511500 667204
rect 325686 656924 325886 657124
rect 333750 656914 334200 657364
rect 415686 656924 415886 657124
rect 423750 656914 424200 657364
rect 505686 656924 505886 657124
rect 513750 656914 514200 657364
rect 55884 655000 56084 655200
rect 63948 654990 64398 655440
rect 145884 655000 146084 655200
rect 153948 654990 154398 655440
rect 235884 655000 236084 655200
rect 243948 654990 244398 655440
rect 57258 646140 57918 646920
rect 60978 646140 61638 646920
rect 147258 646140 147918 646920
rect 150978 646140 151638 646920
rect 237258 646140 237918 646920
rect 327060 648064 327720 648844
rect 330780 648064 331440 648844
rect 417060 648064 417720 648844
rect 420780 648064 421440 648844
rect 507060 648064 507720 648844
rect 510780 648064 511440 648844
rect 240978 646140 241638 646920
rect 417120 591424 417780 592204
rect 57318 589500 57978 590280
rect 61038 589500 61698 590280
rect 147318 589500 147978 590280
rect 151038 589500 151698 590280
rect 237318 589500 237978 590280
rect 241038 589500 241698 590280
rect 327318 589500 327978 590280
rect 331038 589500 331698 590280
rect 420840 591424 421500 592204
rect 507120 591424 507780 592204
rect 510840 591424 511500 592204
rect 415686 581924 415886 582124
rect 423750 581914 424200 582364
rect 505686 581924 505886 582124
rect 513750 581914 514200 582364
rect 55884 580000 56084 580200
rect 63948 579990 64398 580440
rect 145884 580000 146084 580200
rect 153948 579990 154398 580440
rect 235884 580000 236084 580200
rect 243948 579990 244398 580440
rect 325884 580000 326084 580200
rect 333948 579990 334398 580440
rect 57258 571140 57918 571920
rect 60978 571140 61638 571920
rect 147258 571140 147918 571920
rect 150978 571140 151638 571920
rect 237258 571140 237918 571920
rect 240978 571140 241638 571920
rect 327258 571140 327918 571920
rect 417060 573064 417720 573844
rect 420780 573064 421440 573844
rect 507060 573064 507720 573844
rect 510780 573064 511440 573844
rect 330978 571140 331638 571920
rect 64750 508500 65426 509424
rect 154750 508500 155426 509424
rect 244750 508500 245426 509424
rect 334750 508500 335426 509424
rect 424750 508500 425426 509424
rect 514750 508500 515426 509424
rect 57318 500600 57978 501380
rect 61038 500600 61698 501380
rect 147318 500600 147978 501380
rect 151038 500600 151698 501380
rect 237318 500600 237978 501380
rect 241038 500600 241698 501380
rect 327318 500600 327978 501380
rect 331038 500600 331698 501380
rect 417318 500600 417978 501380
rect 421038 500600 421698 501380
rect 507318 500600 507978 501380
rect 511038 500600 511698 501380
rect 229051 493495 229999 494443
rect 320275 492028 320601 492354
rect 55884 491100 56084 491300
rect 63948 491090 64398 491540
rect 340369 491278 340791 491700
rect 415884 491100 416084 491300
rect 423948 491090 424398 491540
rect 505884 491100 506084 491300
rect 513948 491090 514398 491540
rect 139663 486715 140753 487805
rect 158318 486540 159188 487410
rect 249825 486588 251326 488089
rect 57258 482240 57918 483020
rect 60978 482240 61638 483020
rect 147258 482240 147918 483020
rect 150978 482240 151638 483020
rect 237258 482240 237918 483020
rect 240978 482240 241638 483020
rect 327258 482240 327918 483020
rect 330978 482240 331638 483020
rect 417258 482240 417918 483020
rect 420978 482240 421638 483020
rect 507258 482240 507918 483020
rect 510978 482240 511638 483020
rect 52604 474174 53280 475098
rect 142604 474174 143280 475098
rect 232604 474174 233280 475098
rect 322604 474174 323280 475098
rect 412604 474174 413280 475098
rect 502604 474174 503280 475098
rect 64750 388500 65426 389424
rect 154750 388500 155426 389424
rect 244750 388500 245426 389424
rect 334750 388500 335426 389424
rect 424750 388500 425426 389424
rect 514750 388500 515426 389424
rect 57318 380600 57978 381380
rect 61038 380600 61698 381380
rect 147318 380600 147978 381380
rect 151038 380600 151698 381380
rect 237318 380600 237978 381380
rect 241038 380600 241698 381380
rect 327318 380600 327978 381380
rect 331038 380600 331698 381380
rect 417318 380600 417978 381380
rect 421038 380600 421698 381380
rect 507318 380600 507978 381380
rect 511038 380600 511698 381380
rect 229051 373495 229999 374443
rect 320275 372028 320601 372354
rect 340369 371278 340791 371700
rect 415884 371100 416084 371300
rect 423948 371090 424398 371540
rect 505884 371100 506084 371300
rect 513948 371090 514398 371540
rect 49663 366715 50753 367805
rect 68318 366540 69188 367410
rect 139663 366715 140753 367805
rect 158318 366540 159188 367410
rect 249825 366588 251326 368089
rect 57258 362240 57918 363020
rect 60978 362240 61638 363020
rect 147258 362240 147918 363020
rect 150978 362240 151638 363020
rect 237258 362240 237918 363020
rect 240978 362240 241638 363020
rect 327258 362240 327918 363020
rect 330978 362240 331638 363020
rect 417258 362240 417918 363020
rect 420978 362240 421638 363020
rect 507258 362240 507918 363020
rect 510978 362240 511638 363020
rect 52604 354174 53280 355098
rect 142604 354174 143280 355098
rect 232604 354174 233280 355098
rect 322604 354174 323280 355098
rect 412604 354174 413280 355098
rect 502604 354174 503280 355098
rect 64750 268500 65426 269424
rect 153874 268296 154550 269220
rect 245128 268108 245804 269032
rect 334750 268500 335426 269424
rect 424750 268500 425426 269424
rect 514750 268500 515426 269424
rect 57318 260600 57978 261380
rect 61038 260600 61698 261380
rect 146442 260396 147102 261176
rect 150162 260396 150822 261176
rect 237696 260208 238356 260988
rect 241416 260208 242076 260988
rect 327318 260600 327978 261380
rect 331038 260600 331698 261380
rect 417318 260600 417978 261380
rect 421038 260600 421698 261380
rect 507318 260600 507978 261380
rect 511038 260600 511698 261380
rect 319051 253495 319999 254443
rect 55884 251100 56084 251300
rect 63948 251090 64398 251540
rect 230653 251636 230979 251962
rect 145008 250896 145208 251096
rect 153072 250886 153522 251336
rect 250747 250886 251169 251308
rect 339825 246588 341326 248089
rect 409663 246715 410753 247805
rect 428318 246540 429188 247410
rect 499663 246715 500753 247805
rect 518318 246540 519188 247410
rect 57258 242240 57918 243020
rect 60978 242240 61638 243020
rect 146382 242036 147042 242816
rect 150102 242036 150762 242816
rect 237636 241848 238296 242628
rect 241356 241848 242016 242628
rect 327258 242240 327918 243020
rect 330978 242240 331638 243020
rect 417258 242240 417918 243020
rect 420978 242240 421638 243020
rect 507258 242240 507918 243020
rect 510978 242240 511638 243020
rect 52604 234174 53280 235098
rect 141728 233970 142404 234894
rect 232982 233782 233658 234706
rect 322604 234174 323280 235098
rect 412604 234174 413280 235098
rect 502604 234174 503280 235098
rect 57318 154500 57978 155280
rect 61038 154500 61698 155280
rect 147318 154500 147978 155280
rect 151038 154500 151698 155280
rect 237318 154500 237978 155280
rect 241038 154500 241698 155280
rect 327318 154500 327978 155280
rect 331038 154500 331698 155280
rect 417318 154500 417978 155280
rect 421038 154500 421698 155280
rect 507318 154500 507978 155280
rect 511038 154500 511698 155280
rect 55884 145000 56084 145200
rect 63948 144990 64398 145440
rect 145884 145000 146084 145200
rect 153948 144990 154398 145440
rect 235884 145000 236084 145200
rect 243948 144990 244398 145440
rect 325884 145000 326084 145200
rect 333948 144990 334398 145440
rect 415884 145000 416084 145200
rect 423948 144990 424398 145440
rect 505884 145000 506084 145200
rect 513948 144990 514398 145440
rect 57258 136140 57918 136920
rect 60978 136140 61638 136920
rect 147258 136140 147918 136920
rect 150978 136140 151638 136920
rect 237258 136140 237918 136920
rect 240978 136140 241638 136920
rect 327258 136140 327918 136920
rect 330978 136140 331638 136920
rect 417258 136140 417918 136920
rect 420978 136140 421638 136920
rect 507258 136140 507918 136920
rect 510978 136140 511638 136920
rect 57318 64500 57978 65280
rect 61038 64500 61698 65280
rect 147318 64500 147978 65280
rect 151038 64500 151698 65280
rect 237318 64500 237978 65280
rect 241038 64500 241698 65280
rect 327318 64500 327978 65280
rect 331038 64500 331698 65280
rect 417318 64500 417978 65280
rect 421038 64500 421698 65280
rect 507318 64500 507978 65280
rect 511038 64500 511698 65280
rect 55884 55000 56084 55200
rect 63948 54990 64398 55440
rect 145884 55000 146084 55200
rect 153948 54990 154398 55440
rect 235884 55000 236084 55200
rect 243948 54990 244398 55440
rect 325884 55000 326084 55200
rect 333948 54990 334398 55440
rect 415884 55000 416084 55200
rect 423948 54990 424398 55440
rect 505884 55000 506084 55200
rect 513948 54990 514398 55440
rect 57258 46140 57918 46920
rect 60978 46140 61638 46920
rect 147258 46140 147918 46920
rect 150978 46140 151638 46920
rect 237258 46140 237918 46920
rect 240978 46140 241638 46920
rect 327258 46140 327918 46920
rect 330978 46140 331638 46920
rect 417258 46140 417918 46920
rect 420978 46140 421638 46920
rect 507258 46140 507918 46920
rect 510978 46140 511638 46920
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 326940 670624 327900 670864
rect 326940 670144 327060 670624
rect 327780 670144 327900 670624
rect 57138 668700 58098 668940
rect 57138 668220 57258 668700
rect 57978 668220 58098 668700
rect 57138 665280 58098 668220
rect 57138 664500 57318 665280
rect 57978 664500 58098 665280
rect 57138 664140 58098 664500
rect 60858 668700 61818 668940
rect 60858 668220 60978 668700
rect 61698 668220 61818 668700
rect 60858 665280 61818 668220
rect 60858 664500 61038 665280
rect 61698 664500 61818 665280
rect 60858 664140 61818 664500
rect 147138 668700 148098 668940
rect 147138 668220 147258 668700
rect 147978 668220 148098 668700
rect 147138 665280 148098 668220
rect 147138 664500 147318 665280
rect 147978 664500 148098 665280
rect 147138 664140 148098 664500
rect 150858 668700 151818 668940
rect 150858 668220 150978 668700
rect 151698 668220 151818 668700
rect 150858 665280 151818 668220
rect 150858 664500 151038 665280
rect 151698 664500 151818 665280
rect 150858 664140 151818 664500
rect 237138 668700 238098 668940
rect 237138 668220 237258 668700
rect 237978 668220 238098 668700
rect 237138 665280 238098 668220
rect 237138 664500 237318 665280
rect 237978 664500 238098 665280
rect 237138 664140 238098 664500
rect 240858 668700 241818 668940
rect 240858 668220 240978 668700
rect 241698 668220 241818 668700
rect 240858 665280 241818 668220
rect 326940 667204 327900 670144
rect 326940 666424 327120 667204
rect 327780 666424 327900 667204
rect 326940 666064 327900 666424
rect 330660 670624 331620 670864
rect 330660 670144 330780 670624
rect 331500 670144 331620 670624
rect 330660 667204 331620 670144
rect 330660 666424 330840 667204
rect 331500 666424 331620 667204
rect 330660 666064 331620 666424
rect 416940 670624 417900 670864
rect 416940 670144 417060 670624
rect 417780 670144 417900 670624
rect 416940 667204 417900 670144
rect 416940 666424 417120 667204
rect 417780 666424 417900 667204
rect 416940 666064 417900 666424
rect 420660 670624 421620 670864
rect 420660 670144 420780 670624
rect 421500 670144 421620 670624
rect 420660 667204 421620 670144
rect 420660 666424 420840 667204
rect 421500 666424 421620 667204
rect 420660 666064 421620 666424
rect 506940 670624 507900 670864
rect 506940 670144 507060 670624
rect 507780 670144 507900 670624
rect 506940 667204 507900 670144
rect 506940 666424 507120 667204
rect 507780 666424 507900 667204
rect 506940 666064 507900 666424
rect 510660 670624 511620 670864
rect 510660 670144 510780 670624
rect 511500 670144 511620 670624
rect 510660 667204 511620 670144
rect 510660 666424 510840 667204
rect 511500 666424 511620 667204
rect 510660 666064 511620 666424
rect 240858 664500 241038 665280
rect 241698 664500 241818 665280
rect 240858 664140 241818 664500
rect 322962 657184 325924 657882
rect 322962 656864 322996 657184
rect 323316 657124 325924 657184
rect 323316 656924 325686 657124
rect 325886 656924 325924 657124
rect 323316 656864 325924 656924
rect 322962 656556 325924 656864
rect 333544 657779 337084 657864
rect 333544 657648 337093 657779
rect 333544 657364 336368 657648
rect 333544 656914 333750 657364
rect 334200 657014 336368 657364
rect 337020 657014 337093 657648
rect 334200 656914 337093 657014
rect 333544 656903 337093 656914
rect 412962 657184 415924 657882
rect 333544 656594 337084 656903
rect 412962 656864 412996 657184
rect 413316 657124 415924 657184
rect 413316 656924 415686 657124
rect 415886 656924 415924 657124
rect 413316 656864 415924 656924
rect 412962 656556 415924 656864
rect 423544 657779 427084 657864
rect 423544 657648 427093 657779
rect 423544 657364 426368 657648
rect 423544 656914 423750 657364
rect 424200 657014 426368 657364
rect 427020 657014 427093 657648
rect 424200 656914 427093 657014
rect 423544 656903 427093 656914
rect 502962 657184 505924 657882
rect 423544 656594 427084 656903
rect 502962 656864 502996 657184
rect 503316 657124 505924 657184
rect 503316 656924 505686 657124
rect 505886 656924 505924 657124
rect 503316 656864 505924 656924
rect 502962 656556 505924 656864
rect 513544 657779 517084 657864
rect 513544 657648 517093 657779
rect 513544 657364 516368 657648
rect 513544 656914 513750 657364
rect 514200 657014 516368 657364
rect 517020 657014 517093 657648
rect 514200 656914 517093 657014
rect 513544 656903 517093 656914
rect 513544 656594 517084 656903
rect 53160 655260 56122 655958
rect 53160 654940 53194 655260
rect 53514 655200 56122 655260
rect 53514 655000 55884 655200
rect 56084 655000 56122 655200
rect 53514 654940 56122 655000
rect 53160 654632 56122 654940
rect 63742 655855 67282 655940
rect 63742 655724 67291 655855
rect 63742 655440 66566 655724
rect 63742 654990 63948 655440
rect 64398 655090 66566 655440
rect 67218 655090 67291 655724
rect 64398 654990 67291 655090
rect 63742 654979 67291 654990
rect 143160 655260 146122 655958
rect 63742 654670 67282 654979
rect 143160 654940 143194 655260
rect 143514 655200 146122 655260
rect 143514 655000 145884 655200
rect 146084 655000 146122 655200
rect 143514 654940 146122 655000
rect 143160 654632 146122 654940
rect 153742 655855 157282 655940
rect 153742 655724 157291 655855
rect 153742 655440 156566 655724
rect 153742 654990 153948 655440
rect 154398 655090 156566 655440
rect 157218 655090 157291 655724
rect 154398 654990 157291 655090
rect 153742 654979 157291 654990
rect 233160 655260 236122 655958
rect 153742 654670 157282 654979
rect 233160 654940 233194 655260
rect 233514 655200 236122 655260
rect 233514 655000 235884 655200
rect 236084 655000 236122 655200
rect 233514 654940 236122 655000
rect 233160 654632 236122 654940
rect 243742 655855 247282 655940
rect 243742 655724 247291 655855
rect 243742 655440 246566 655724
rect 243742 654990 243948 655440
rect 244398 655090 246566 655440
rect 247218 655090 247291 655724
rect 244398 654990 247291 655090
rect 243742 654979 247291 654990
rect 243742 654670 247282 654979
rect 326880 648844 327840 649204
rect 326880 648064 327060 648844
rect 327720 648064 327840 648844
rect 57078 646920 58038 647280
rect 57078 646140 57258 646920
rect 57918 646140 58038 646920
rect 57078 643200 58038 646140
rect 57078 642720 57198 643200
rect 57918 642720 58038 643200
rect 57078 642480 58038 642720
rect 60798 646920 61758 647280
rect 60798 646140 60978 646920
rect 61638 646140 61758 646920
rect 60798 643200 61758 646140
rect 60798 642720 60918 643200
rect 61638 642720 61758 643200
rect 60798 642480 61758 642720
rect 147078 646920 148038 647280
rect 147078 646140 147258 646920
rect 147918 646140 148038 646920
rect 147078 643200 148038 646140
rect 147078 642720 147198 643200
rect 147918 642720 148038 643200
rect 147078 642480 148038 642720
rect 150798 646920 151758 647280
rect 150798 646140 150978 646920
rect 151638 646140 151758 646920
rect 150798 643200 151758 646140
rect 150798 642720 150918 643200
rect 151638 642720 151758 643200
rect 150798 642480 151758 642720
rect 237078 646920 238038 647280
rect 237078 646140 237258 646920
rect 237918 646140 238038 646920
rect 237078 643200 238038 646140
rect 237078 642720 237198 643200
rect 237918 642720 238038 643200
rect 237078 642480 238038 642720
rect 240798 646920 241758 647280
rect 240798 646140 240978 646920
rect 241638 646140 241758 646920
rect 240798 643200 241758 646140
rect 326880 645124 327840 648064
rect 326880 644644 327000 645124
rect 327720 644644 327840 645124
rect 326880 644404 327840 644644
rect 330600 648844 331560 649204
rect 330600 648064 330780 648844
rect 331440 648064 331560 648844
rect 330600 645124 331560 648064
rect 330600 644644 330720 645124
rect 331440 644644 331560 645124
rect 330600 644404 331560 644644
rect 416880 648844 417840 649204
rect 416880 648064 417060 648844
rect 417720 648064 417840 648844
rect 416880 645124 417840 648064
rect 416880 644644 417000 645124
rect 417720 644644 417840 645124
rect 416880 644404 417840 644644
rect 420600 648844 421560 649204
rect 420600 648064 420780 648844
rect 421440 648064 421560 648844
rect 420600 645124 421560 648064
rect 420600 644644 420720 645124
rect 421440 644644 421560 645124
rect 420600 644404 421560 644644
rect 506880 648844 507840 649204
rect 506880 648064 507060 648844
rect 507720 648064 507840 648844
rect 506880 645124 507840 648064
rect 506880 644644 507000 645124
rect 507720 644644 507840 645124
rect 506880 644404 507840 644644
rect 510600 648844 511560 649204
rect 510600 648064 510780 648844
rect 511440 648064 511560 648844
rect 510600 645124 511560 648064
rect 510600 644644 510720 645124
rect 511440 644644 511560 645124
rect 510600 644404 511560 644644
rect 240798 642720 240918 643200
rect 241638 642720 241758 643200
rect 240798 642480 241758 642720
rect 416940 595624 417900 595864
rect 416940 595144 417060 595624
rect 417780 595144 417900 595624
rect 57138 593700 58098 593940
rect 57138 593220 57258 593700
rect 57978 593220 58098 593700
rect 57138 590280 58098 593220
rect 57138 589500 57318 590280
rect 57978 589500 58098 590280
rect 57138 589140 58098 589500
rect 60858 593700 61818 593940
rect 60858 593220 60978 593700
rect 61698 593220 61818 593700
rect 60858 590280 61818 593220
rect 60858 589500 61038 590280
rect 61698 589500 61818 590280
rect 60858 589140 61818 589500
rect 147138 593700 148098 593940
rect 147138 593220 147258 593700
rect 147978 593220 148098 593700
rect 147138 590280 148098 593220
rect 147138 589500 147318 590280
rect 147978 589500 148098 590280
rect 147138 589140 148098 589500
rect 150858 593700 151818 593940
rect 150858 593220 150978 593700
rect 151698 593220 151818 593700
rect 150858 590280 151818 593220
rect 150858 589500 151038 590280
rect 151698 589500 151818 590280
rect 150858 589140 151818 589500
rect 237138 593700 238098 593940
rect 237138 593220 237258 593700
rect 237978 593220 238098 593700
rect 237138 590280 238098 593220
rect 237138 589500 237318 590280
rect 237978 589500 238098 590280
rect 237138 589140 238098 589500
rect 240858 593700 241818 593940
rect 240858 593220 240978 593700
rect 241698 593220 241818 593700
rect 240858 590280 241818 593220
rect 240858 589500 241038 590280
rect 241698 589500 241818 590280
rect 240858 589140 241818 589500
rect 327138 593700 328098 593940
rect 327138 593220 327258 593700
rect 327978 593220 328098 593700
rect 327138 590280 328098 593220
rect 327138 589500 327318 590280
rect 327978 589500 328098 590280
rect 327138 589140 328098 589500
rect 330858 593700 331818 593940
rect 330858 593220 330978 593700
rect 331698 593220 331818 593700
rect 330858 590280 331818 593220
rect 416940 592204 417900 595144
rect 416940 591424 417120 592204
rect 417780 591424 417900 592204
rect 416940 591064 417900 591424
rect 420660 595624 421620 595864
rect 420660 595144 420780 595624
rect 421500 595144 421620 595624
rect 420660 592204 421620 595144
rect 420660 591424 420840 592204
rect 421500 591424 421620 592204
rect 420660 591064 421620 591424
rect 506940 595624 507900 595864
rect 506940 595144 507060 595624
rect 507780 595144 507900 595624
rect 506940 592204 507900 595144
rect 506940 591424 507120 592204
rect 507780 591424 507900 592204
rect 506940 591064 507900 591424
rect 510660 595624 511620 595864
rect 510660 595144 510780 595624
rect 511500 595144 511620 595624
rect 510660 592204 511620 595144
rect 510660 591424 510840 592204
rect 511500 591424 511620 592204
rect 510660 591064 511620 591424
rect 330858 589500 331038 590280
rect 331698 589500 331818 590280
rect 330858 589140 331818 589500
rect 412962 582184 415924 582882
rect 412962 581864 412996 582184
rect 413316 582124 415924 582184
rect 413316 581924 415686 582124
rect 415886 581924 415924 582124
rect 413316 581864 415924 581924
rect 412962 581556 415924 581864
rect 423544 582779 427084 582864
rect 423544 582648 427093 582779
rect 423544 582364 426368 582648
rect 423544 581914 423750 582364
rect 424200 582014 426368 582364
rect 427020 582014 427093 582648
rect 424200 581914 427093 582014
rect 423544 581903 427093 581914
rect 502962 582184 505924 582882
rect 423544 581594 427084 581903
rect 502962 581864 502996 582184
rect 503316 582124 505924 582184
rect 503316 581924 505686 582124
rect 505886 581924 505924 582124
rect 503316 581864 505924 581924
rect 502962 581556 505924 581864
rect 513544 582779 517084 582864
rect 513544 582648 517093 582779
rect 513544 582364 516368 582648
rect 513544 581914 513750 582364
rect 514200 582014 516368 582364
rect 517020 582014 517093 582648
rect 514200 581914 517093 582014
rect 513544 581903 517093 581914
rect 513544 581594 517084 581903
rect 53160 580260 56122 580958
rect 53160 579940 53194 580260
rect 53514 580200 56122 580260
rect 53514 580000 55884 580200
rect 56084 580000 56122 580200
rect 53514 579940 56122 580000
rect 53160 579632 56122 579940
rect 63742 580855 67282 580940
rect 63742 580724 67291 580855
rect 63742 580440 66566 580724
rect 63742 579990 63948 580440
rect 64398 580090 66566 580440
rect 67218 580090 67291 580724
rect 64398 579990 67291 580090
rect 63742 579979 67291 579990
rect 143160 580260 146122 580958
rect 63742 579670 67282 579979
rect 143160 579940 143194 580260
rect 143514 580200 146122 580260
rect 143514 580000 145884 580200
rect 146084 580000 146122 580200
rect 143514 579940 146122 580000
rect 143160 579632 146122 579940
rect 153742 580855 157282 580940
rect 153742 580724 157291 580855
rect 153742 580440 156566 580724
rect 153742 579990 153948 580440
rect 154398 580090 156566 580440
rect 157218 580090 157291 580724
rect 154398 579990 157291 580090
rect 153742 579979 157291 579990
rect 233160 580260 236122 580958
rect 153742 579670 157282 579979
rect 233160 579940 233194 580260
rect 233514 580200 236122 580260
rect 233514 580000 235884 580200
rect 236084 580000 236122 580200
rect 233514 579940 236122 580000
rect 233160 579632 236122 579940
rect 243742 580855 247282 580940
rect 243742 580724 247291 580855
rect 243742 580440 246566 580724
rect 243742 579990 243948 580440
rect 244398 580090 246566 580440
rect 247218 580090 247291 580724
rect 244398 579990 247291 580090
rect 243742 579979 247291 579990
rect 323160 580260 326122 580958
rect 243742 579670 247282 579979
rect 323160 579940 323194 580260
rect 323514 580200 326122 580260
rect 323514 580000 325884 580200
rect 326084 580000 326122 580200
rect 323514 579940 326122 580000
rect 323160 579632 326122 579940
rect 333742 580855 337282 580940
rect 333742 580724 337291 580855
rect 333742 580440 336566 580724
rect 333742 579990 333948 580440
rect 334398 580090 336566 580440
rect 337218 580090 337291 580724
rect 334398 579990 337291 580090
rect 333742 579979 337291 579990
rect 333742 579670 337282 579979
rect 416880 573844 417840 574204
rect 416880 573064 417060 573844
rect 417720 573064 417840 573844
rect 57078 571920 58038 572280
rect 57078 571140 57258 571920
rect 57918 571140 58038 571920
rect 57078 568200 58038 571140
rect 57078 567720 57198 568200
rect 57918 567720 58038 568200
rect 57078 567480 58038 567720
rect 60798 571920 61758 572280
rect 60798 571140 60978 571920
rect 61638 571140 61758 571920
rect 60798 568200 61758 571140
rect 60798 567720 60918 568200
rect 61638 567720 61758 568200
rect 60798 567480 61758 567720
rect 147078 571920 148038 572280
rect 147078 571140 147258 571920
rect 147918 571140 148038 571920
rect 147078 568200 148038 571140
rect 147078 567720 147198 568200
rect 147918 567720 148038 568200
rect 147078 567480 148038 567720
rect 150798 571920 151758 572280
rect 150798 571140 150978 571920
rect 151638 571140 151758 571920
rect 150798 568200 151758 571140
rect 150798 567720 150918 568200
rect 151638 567720 151758 568200
rect 150798 567480 151758 567720
rect 237078 571920 238038 572280
rect 237078 571140 237258 571920
rect 237918 571140 238038 571920
rect 237078 568200 238038 571140
rect 237078 567720 237198 568200
rect 237918 567720 238038 568200
rect 237078 567480 238038 567720
rect 240798 571920 241758 572280
rect 240798 571140 240978 571920
rect 241638 571140 241758 571920
rect 240798 568200 241758 571140
rect 240798 567720 240918 568200
rect 241638 567720 241758 568200
rect 240798 567480 241758 567720
rect 327078 571920 328038 572280
rect 327078 571140 327258 571920
rect 327918 571140 328038 571920
rect 327078 568200 328038 571140
rect 327078 567720 327198 568200
rect 327918 567720 328038 568200
rect 327078 567480 328038 567720
rect 330798 571920 331758 572280
rect 330798 571140 330978 571920
rect 331638 571140 331758 571920
rect 330798 568200 331758 571140
rect 416880 570124 417840 573064
rect 416880 569644 417000 570124
rect 417720 569644 417840 570124
rect 416880 569404 417840 569644
rect 420600 573844 421560 574204
rect 420600 573064 420780 573844
rect 421440 573064 421560 573844
rect 420600 570124 421560 573064
rect 420600 569644 420720 570124
rect 421440 569644 421560 570124
rect 420600 569404 421560 569644
rect 506880 573844 507840 574204
rect 506880 573064 507060 573844
rect 507720 573064 507840 573844
rect 506880 570124 507840 573064
rect 506880 569644 507000 570124
rect 507720 569644 507840 570124
rect 506880 569404 507840 569644
rect 510600 573844 511560 574204
rect 510600 573064 510780 573844
rect 511440 573064 511560 573844
rect 510600 570124 511560 573064
rect 510600 569644 510720 570124
rect 511440 569644 511560 570124
rect 510600 569404 511560 569644
rect 330798 567720 330918 568200
rect 331638 567720 331758 568200
rect 330798 567480 331758 567720
rect 63816 516794 66396 517438
rect 63816 515116 64332 516794
rect 65752 515116 66396 516794
rect 63816 509424 66396 515116
rect 63816 508500 64750 509424
rect 65426 508500 66396 509424
rect 63816 507892 66396 508500
rect 153816 516794 156396 517438
rect 153816 515116 154332 516794
rect 155752 515116 156396 516794
rect 153816 509424 156396 515116
rect 153816 508500 154750 509424
rect 155426 508500 156396 509424
rect 153816 507892 156396 508500
rect 243816 516794 246396 517438
rect 243816 515116 244332 516794
rect 245752 515116 246396 516794
rect 243816 509424 246396 515116
rect 243816 508500 244750 509424
rect 245426 508500 246396 509424
rect 243816 507892 246396 508500
rect 333816 516794 336396 517438
rect 333816 515116 334332 516794
rect 335752 515116 336396 516794
rect 333816 509424 336396 515116
rect 333816 508500 334750 509424
rect 335426 508500 336396 509424
rect 333816 507892 336396 508500
rect 423816 516794 426396 517438
rect 423816 515116 424332 516794
rect 425752 515116 426396 516794
rect 423816 509424 426396 515116
rect 423816 508500 424750 509424
rect 425426 508500 426396 509424
rect 423816 507892 426396 508500
rect 513816 516794 516396 517438
rect 513816 515116 514332 516794
rect 515752 515116 516396 516794
rect 513816 509424 516396 515116
rect 513816 508500 514750 509424
rect 515426 508500 516396 509424
rect 513816 507892 516396 508500
rect 57138 504800 58098 505040
rect 57138 504320 57258 504800
rect 57978 504320 58098 504800
rect 57138 501380 58098 504320
rect 57138 500600 57318 501380
rect 57978 500600 58098 501380
rect 57138 500240 58098 500600
rect 60858 504800 61818 505040
rect 60858 504320 60978 504800
rect 61698 504320 61818 504800
rect 60858 501380 61818 504320
rect 60858 500600 61038 501380
rect 61698 500600 61818 501380
rect 60858 500240 61818 500600
rect 147138 504800 148098 505040
rect 147138 504320 147258 504800
rect 147978 504320 148098 504800
rect 147138 501380 148098 504320
rect 147138 500600 147318 501380
rect 147978 500600 148098 501380
rect 147138 500240 148098 500600
rect 150858 504800 151818 505040
rect 150858 504320 150978 504800
rect 151698 504320 151818 504800
rect 150858 501380 151818 504320
rect 150858 500600 151038 501380
rect 151698 500600 151818 501380
rect 150858 500240 151818 500600
rect 237138 504800 238098 505040
rect 237138 504320 237258 504800
rect 237978 504320 238098 504800
rect 237138 501380 238098 504320
rect 237138 500600 237318 501380
rect 237978 500600 238098 501380
rect 237138 500240 238098 500600
rect 240858 504800 241818 505040
rect 240858 504320 240978 504800
rect 241698 504320 241818 504800
rect 240858 501380 241818 504320
rect 240858 500600 241038 501380
rect 241698 500600 241818 501380
rect 240858 500240 241818 500600
rect 327138 504800 328098 505040
rect 327138 504320 327258 504800
rect 327978 504320 328098 504800
rect 327138 501380 328098 504320
rect 327138 500600 327318 501380
rect 327978 500600 328098 501380
rect 327138 500240 328098 500600
rect 330858 504800 331818 505040
rect 330858 504320 330978 504800
rect 331698 504320 331818 504800
rect 330858 501380 331818 504320
rect 330858 500600 331038 501380
rect 331698 500600 331818 501380
rect 330858 500240 331818 500600
rect 417138 504800 418098 505040
rect 417138 504320 417258 504800
rect 417978 504320 418098 504800
rect 417138 501380 418098 504320
rect 417138 500600 417318 501380
rect 417978 500600 418098 501380
rect 417138 500240 418098 500600
rect 420858 504800 421818 505040
rect 420858 504320 420978 504800
rect 421698 504320 421818 504800
rect 420858 501380 421818 504320
rect 420858 500600 421038 501380
rect 421698 500600 421818 501380
rect 420858 500240 421818 500600
rect 507138 504800 508098 505040
rect 507138 504320 507258 504800
rect 507978 504320 508098 504800
rect 507138 501380 508098 504320
rect 507138 500600 507318 501380
rect 507978 500600 508098 501380
rect 507138 500240 508098 500600
rect 510858 504800 511818 505040
rect 510858 504320 510978 504800
rect 511698 504320 511818 504800
rect 510858 501380 511818 504320
rect 510858 500600 511038 501380
rect 511698 500600 511818 501380
rect 510858 500240 511818 500600
rect 229050 494443 230000 494444
rect 227669 493495 229051 494443
rect 229999 493495 230000 494443
rect 53160 491360 56122 492058
rect 53160 491040 53194 491360
rect 53514 491300 56122 491360
rect 53514 491100 55884 491300
rect 56084 491100 56122 491300
rect 53514 491040 56122 491100
rect 53160 490732 56122 491040
rect 63742 491955 67282 492040
rect 63742 491824 67291 491955
rect 63742 491540 66566 491824
rect 63742 491090 63948 491540
rect 64398 491190 66566 491540
rect 67218 491190 67291 491824
rect 64398 491090 67291 491190
rect 63742 491079 67291 491090
rect 227669 491774 228617 493495
rect 229050 493494 230000 493495
rect 320274 492354 320602 492355
rect 63742 490770 67282 491079
rect 319627 492028 320275 492354
rect 320601 492028 320602 492354
rect 319627 491749 319953 492028
rect 320274 492027 320602 492028
rect 340368 491700 340792 491701
rect 340368 491278 340369 491700
rect 340791 491278 341405 491700
rect 413160 491360 416122 492058
rect 340368 491277 340792 491278
rect 413160 491040 413194 491360
rect 413514 491300 416122 491360
rect 413514 491100 415884 491300
rect 416084 491100 416122 491300
rect 413514 491040 416122 491100
rect 413160 490732 416122 491040
rect 423742 491955 427282 492040
rect 423742 491824 427291 491955
rect 423742 491540 426566 491824
rect 423742 491090 423948 491540
rect 424398 491190 426566 491540
rect 427218 491190 427291 491824
rect 424398 491090 427291 491190
rect 423742 491079 427291 491090
rect 503160 491360 506122 492058
rect 423742 490770 427282 491079
rect 503160 491040 503194 491360
rect 503514 491300 506122 491360
rect 503514 491100 505884 491300
rect 506084 491100 506122 491300
rect 503514 491040 506122 491100
rect 503160 490732 506122 491040
rect 513742 491955 517282 492040
rect 513742 491824 517291 491955
rect 513742 491540 516566 491824
rect 513742 491090 513948 491540
rect 514398 491190 516566 491540
rect 517218 491190 517291 491824
rect 514398 491090 517291 491190
rect 513742 491079 517291 491090
rect 513742 490770 517282 491079
rect 249825 488090 251326 490662
rect 249824 488089 251327 488090
rect 139662 487805 140754 487806
rect 139662 486715 139663 487805
rect 140753 486715 140754 487805
rect 139662 486714 140754 486715
rect 158317 487410 159189 487411
rect 139663 485900 140753 486714
rect 158317 486540 158318 487410
rect 159188 486540 160183 487410
rect 249824 486588 249825 488089
rect 251326 486588 251327 488089
rect 249824 486587 251327 486588
rect 158317 486539 159189 486540
rect 57078 483020 58038 483380
rect 57078 482240 57258 483020
rect 57918 482240 58038 483020
rect 57078 479300 58038 482240
rect 57078 478820 57198 479300
rect 57918 478820 58038 479300
rect 57078 478580 58038 478820
rect 60798 483020 61758 483380
rect 60798 482240 60978 483020
rect 61638 482240 61758 483020
rect 60798 479300 61758 482240
rect 60798 478820 60918 479300
rect 61638 478820 61758 479300
rect 60798 478580 61758 478820
rect 147078 483020 148038 483380
rect 147078 482240 147258 483020
rect 147918 482240 148038 483020
rect 147078 479300 148038 482240
rect 147078 478820 147198 479300
rect 147918 478820 148038 479300
rect 147078 478580 148038 478820
rect 150798 483020 151758 483380
rect 150798 482240 150978 483020
rect 151638 482240 151758 483020
rect 150798 479300 151758 482240
rect 150798 478820 150918 479300
rect 151638 478820 151758 479300
rect 150798 478580 151758 478820
rect 237078 483020 238038 483380
rect 237078 482240 237258 483020
rect 237918 482240 238038 483020
rect 237078 479300 238038 482240
rect 237078 478820 237198 479300
rect 237918 478820 238038 479300
rect 237078 478580 238038 478820
rect 240798 483020 241758 483380
rect 240798 482240 240978 483020
rect 241638 482240 241758 483020
rect 240798 479300 241758 482240
rect 240798 478820 240918 479300
rect 241638 478820 241758 479300
rect 240798 478580 241758 478820
rect 327078 483020 328038 483380
rect 327078 482240 327258 483020
rect 327918 482240 328038 483020
rect 327078 479300 328038 482240
rect 327078 478820 327198 479300
rect 327918 478820 328038 479300
rect 327078 478580 328038 478820
rect 330798 483020 331758 483380
rect 330798 482240 330978 483020
rect 331638 482240 331758 483020
rect 330798 479300 331758 482240
rect 330798 478820 330918 479300
rect 331638 478820 331758 479300
rect 330798 478580 331758 478820
rect 417078 483020 418038 483380
rect 417078 482240 417258 483020
rect 417918 482240 418038 483020
rect 417078 479300 418038 482240
rect 417078 478820 417198 479300
rect 417918 478820 418038 479300
rect 417078 478580 418038 478820
rect 420798 483020 421758 483380
rect 420798 482240 420978 483020
rect 421638 482240 421758 483020
rect 420798 479300 421758 482240
rect 420798 478820 420918 479300
rect 421638 478820 421758 479300
rect 420798 478580 421758 478820
rect 507078 483020 508038 483380
rect 507078 482240 507258 483020
rect 507918 482240 508038 483020
rect 507078 479300 508038 482240
rect 507078 478820 507198 479300
rect 507918 478820 508038 479300
rect 507078 478580 508038 478820
rect 510798 483020 511758 483380
rect 510798 482240 510978 483020
rect 511638 482240 511758 483020
rect 510798 479300 511758 482240
rect 510798 478820 510918 479300
rect 511638 478820 511758 479300
rect 510798 478580 511758 478820
rect 51754 475098 54334 475446
rect 51754 474174 52604 475098
rect 53280 474174 54334 475098
rect 51754 468222 54334 474174
rect 51754 466544 52334 468222
rect 53754 466544 54334 468222
rect 51754 465900 54334 466544
rect 141754 475098 144334 475446
rect 141754 474174 142604 475098
rect 143280 474174 144334 475098
rect 141754 468222 144334 474174
rect 141754 466544 142334 468222
rect 143754 466544 144334 468222
rect 141754 465900 144334 466544
rect 231754 475098 234334 475446
rect 231754 474174 232604 475098
rect 233280 474174 234334 475098
rect 231754 468222 234334 474174
rect 231754 466544 232334 468222
rect 233754 466544 234334 468222
rect 231754 465900 234334 466544
rect 321754 475098 324334 475446
rect 321754 474174 322604 475098
rect 323280 474174 324334 475098
rect 321754 468222 324334 474174
rect 321754 466544 322334 468222
rect 323754 466544 324334 468222
rect 321754 465900 324334 466544
rect 411754 475098 414334 475446
rect 411754 474174 412604 475098
rect 413280 474174 414334 475098
rect 411754 468222 414334 474174
rect 411754 466544 412334 468222
rect 413754 466544 414334 468222
rect 411754 465900 414334 466544
rect 501754 475098 504334 475446
rect 501754 474174 502604 475098
rect 503280 474174 504334 475098
rect 501754 468222 504334 474174
rect 501754 466544 502334 468222
rect 503754 466544 504334 468222
rect 501754 465900 504334 466544
rect 63816 396794 66396 397438
rect 63816 395116 64332 396794
rect 65752 395116 66396 396794
rect 63816 389424 66396 395116
rect 63816 388500 64750 389424
rect 65426 388500 66396 389424
rect 63816 387892 66396 388500
rect 153816 396794 156396 397438
rect 153816 395116 154332 396794
rect 155752 395116 156396 396794
rect 153816 389424 156396 395116
rect 153816 388500 154750 389424
rect 155426 388500 156396 389424
rect 153816 387892 156396 388500
rect 243816 396794 246396 397438
rect 243816 395116 244332 396794
rect 245752 395116 246396 396794
rect 243816 389424 246396 395116
rect 243816 388500 244750 389424
rect 245426 388500 246396 389424
rect 243816 387892 246396 388500
rect 333816 396794 336396 397438
rect 333816 395116 334332 396794
rect 335752 395116 336396 396794
rect 333816 389424 336396 395116
rect 333816 388500 334750 389424
rect 335426 388500 336396 389424
rect 333816 387892 336396 388500
rect 423816 396794 426396 397438
rect 423816 395116 424332 396794
rect 425752 395116 426396 396794
rect 423816 389424 426396 395116
rect 423816 388500 424750 389424
rect 425426 388500 426396 389424
rect 423816 387892 426396 388500
rect 513816 396794 516396 397438
rect 513816 395116 514332 396794
rect 515752 395116 516396 396794
rect 513816 389424 516396 395116
rect 513816 388500 514750 389424
rect 515426 388500 516396 389424
rect 513816 387892 516396 388500
rect 57138 384800 58098 385040
rect 57138 384320 57258 384800
rect 57978 384320 58098 384800
rect 57138 381380 58098 384320
rect 57138 380600 57318 381380
rect 57978 380600 58098 381380
rect 57138 380240 58098 380600
rect 60858 384800 61818 385040
rect 60858 384320 60978 384800
rect 61698 384320 61818 384800
rect 60858 381380 61818 384320
rect 60858 380600 61038 381380
rect 61698 380600 61818 381380
rect 60858 380240 61818 380600
rect 147138 384800 148098 385040
rect 147138 384320 147258 384800
rect 147978 384320 148098 384800
rect 147138 381380 148098 384320
rect 147138 380600 147318 381380
rect 147978 380600 148098 381380
rect 147138 380240 148098 380600
rect 150858 384800 151818 385040
rect 150858 384320 150978 384800
rect 151698 384320 151818 384800
rect 150858 381380 151818 384320
rect 150858 380600 151038 381380
rect 151698 380600 151818 381380
rect 150858 380240 151818 380600
rect 237138 384800 238098 385040
rect 237138 384320 237258 384800
rect 237978 384320 238098 384800
rect 237138 381380 238098 384320
rect 237138 380600 237318 381380
rect 237978 380600 238098 381380
rect 237138 380240 238098 380600
rect 240858 384800 241818 385040
rect 240858 384320 240978 384800
rect 241698 384320 241818 384800
rect 240858 381380 241818 384320
rect 240858 380600 241038 381380
rect 241698 380600 241818 381380
rect 240858 380240 241818 380600
rect 327138 384800 328098 385040
rect 327138 384320 327258 384800
rect 327978 384320 328098 384800
rect 327138 381380 328098 384320
rect 327138 380600 327318 381380
rect 327978 380600 328098 381380
rect 327138 380240 328098 380600
rect 330858 384800 331818 385040
rect 330858 384320 330978 384800
rect 331698 384320 331818 384800
rect 330858 381380 331818 384320
rect 330858 380600 331038 381380
rect 331698 380600 331818 381380
rect 330858 380240 331818 380600
rect 417138 384800 418098 385040
rect 417138 384320 417258 384800
rect 417978 384320 418098 384800
rect 417138 381380 418098 384320
rect 417138 380600 417318 381380
rect 417978 380600 418098 381380
rect 417138 380240 418098 380600
rect 420858 384800 421818 385040
rect 420858 384320 420978 384800
rect 421698 384320 421818 384800
rect 420858 381380 421818 384320
rect 420858 380600 421038 381380
rect 421698 380600 421818 381380
rect 420858 380240 421818 380600
rect 507138 384800 508098 385040
rect 507138 384320 507258 384800
rect 507978 384320 508098 384800
rect 507138 381380 508098 384320
rect 507138 380600 507318 381380
rect 507978 380600 508098 381380
rect 507138 380240 508098 380600
rect 510858 384800 511818 385040
rect 510858 384320 510978 384800
rect 511698 384320 511818 384800
rect 510858 381380 511818 384320
rect 510858 380600 511038 381380
rect 511698 380600 511818 381380
rect 510858 380240 511818 380600
rect 229050 374443 230000 374444
rect 227669 373495 229051 374443
rect 229999 373495 230000 374443
rect 227669 371774 228617 373495
rect 229050 373494 230000 373495
rect 320274 372354 320602 372355
rect 319627 372028 320275 372354
rect 320601 372028 320602 372354
rect 319627 371749 319953 372028
rect 320274 372027 320602 372028
rect 340368 371700 340792 371701
rect 340368 371278 340369 371700
rect 340791 371278 341405 371700
rect 413160 371360 416122 372058
rect 340368 371277 340792 371278
rect 413160 371040 413194 371360
rect 413514 371300 416122 371360
rect 413514 371100 415884 371300
rect 416084 371100 416122 371300
rect 413514 371040 416122 371100
rect 413160 370732 416122 371040
rect 423742 371955 427282 372040
rect 423742 371824 427291 371955
rect 423742 371540 426566 371824
rect 423742 371090 423948 371540
rect 424398 371190 426566 371540
rect 427218 371190 427291 371824
rect 424398 371090 427291 371190
rect 423742 371079 427291 371090
rect 503160 371360 506122 372058
rect 423742 370770 427282 371079
rect 503160 371040 503194 371360
rect 503514 371300 506122 371360
rect 503514 371100 505884 371300
rect 506084 371100 506122 371300
rect 503514 371040 506122 371100
rect 503160 370732 506122 371040
rect 513742 371955 517282 372040
rect 513742 371824 517291 371955
rect 513742 371540 516566 371824
rect 513742 371090 513948 371540
rect 514398 371190 516566 371540
rect 517218 371190 517291 371824
rect 514398 371090 517291 371190
rect 513742 371079 517291 371090
rect 513742 370770 517282 371079
rect 249825 368090 251326 370662
rect 249824 368089 251327 368090
rect 49662 367805 50754 367806
rect 49662 366715 49663 367805
rect 50753 366715 50754 367805
rect 139662 367805 140754 367806
rect 49662 366714 50754 366715
rect 68317 367410 69189 367411
rect 49663 365900 50753 366714
rect 68317 366540 68318 367410
rect 69188 366540 70183 367410
rect 139662 366715 139663 367805
rect 140753 366715 140754 367805
rect 139662 366714 140754 366715
rect 158317 367410 159189 367411
rect 68317 366539 69189 366540
rect 139663 365900 140753 366714
rect 158317 366540 158318 367410
rect 159188 366540 160183 367410
rect 249824 366588 249825 368089
rect 251326 366588 251327 368089
rect 249824 366587 251327 366588
rect 158317 366539 159189 366540
rect 57078 363020 58038 363380
rect 57078 362240 57258 363020
rect 57918 362240 58038 363020
rect 57078 359300 58038 362240
rect 57078 358820 57198 359300
rect 57918 358820 58038 359300
rect 57078 358580 58038 358820
rect 60798 363020 61758 363380
rect 60798 362240 60978 363020
rect 61638 362240 61758 363020
rect 60798 359300 61758 362240
rect 60798 358820 60918 359300
rect 61638 358820 61758 359300
rect 60798 358580 61758 358820
rect 147078 363020 148038 363380
rect 147078 362240 147258 363020
rect 147918 362240 148038 363020
rect 147078 359300 148038 362240
rect 147078 358820 147198 359300
rect 147918 358820 148038 359300
rect 147078 358580 148038 358820
rect 150798 363020 151758 363380
rect 150798 362240 150978 363020
rect 151638 362240 151758 363020
rect 150798 359300 151758 362240
rect 150798 358820 150918 359300
rect 151638 358820 151758 359300
rect 150798 358580 151758 358820
rect 237078 363020 238038 363380
rect 237078 362240 237258 363020
rect 237918 362240 238038 363020
rect 237078 359300 238038 362240
rect 237078 358820 237198 359300
rect 237918 358820 238038 359300
rect 237078 358580 238038 358820
rect 240798 363020 241758 363380
rect 240798 362240 240978 363020
rect 241638 362240 241758 363020
rect 240798 359300 241758 362240
rect 240798 358820 240918 359300
rect 241638 358820 241758 359300
rect 240798 358580 241758 358820
rect 327078 363020 328038 363380
rect 327078 362240 327258 363020
rect 327918 362240 328038 363020
rect 327078 359300 328038 362240
rect 327078 358820 327198 359300
rect 327918 358820 328038 359300
rect 327078 358580 328038 358820
rect 330798 363020 331758 363380
rect 330798 362240 330978 363020
rect 331638 362240 331758 363020
rect 330798 359300 331758 362240
rect 330798 358820 330918 359300
rect 331638 358820 331758 359300
rect 330798 358580 331758 358820
rect 417078 363020 418038 363380
rect 417078 362240 417258 363020
rect 417918 362240 418038 363020
rect 417078 359300 418038 362240
rect 417078 358820 417198 359300
rect 417918 358820 418038 359300
rect 417078 358580 418038 358820
rect 420798 363020 421758 363380
rect 420798 362240 420978 363020
rect 421638 362240 421758 363020
rect 420798 359300 421758 362240
rect 420798 358820 420918 359300
rect 421638 358820 421758 359300
rect 420798 358580 421758 358820
rect 507078 363020 508038 363380
rect 507078 362240 507258 363020
rect 507918 362240 508038 363020
rect 507078 359300 508038 362240
rect 507078 358820 507198 359300
rect 507918 358820 508038 359300
rect 507078 358580 508038 358820
rect 510798 363020 511758 363380
rect 510798 362240 510978 363020
rect 511638 362240 511758 363020
rect 510798 359300 511758 362240
rect 510798 358820 510918 359300
rect 511638 358820 511758 359300
rect 510798 358580 511758 358820
rect 51754 355098 54334 355446
rect 51754 354174 52604 355098
rect 53280 354174 54334 355098
rect 51754 348222 54334 354174
rect 51754 346544 52334 348222
rect 53754 346544 54334 348222
rect 51754 345900 54334 346544
rect 141754 355098 144334 355446
rect 141754 354174 142604 355098
rect 143280 354174 144334 355098
rect 141754 348222 144334 354174
rect 141754 346544 142334 348222
rect 143754 346544 144334 348222
rect 141754 345900 144334 346544
rect 231754 355098 234334 355446
rect 231754 354174 232604 355098
rect 233280 354174 234334 355098
rect 231754 348222 234334 354174
rect 231754 346544 232334 348222
rect 233754 346544 234334 348222
rect 231754 345900 234334 346544
rect 321754 355098 324334 355446
rect 321754 354174 322604 355098
rect 323280 354174 324334 355098
rect 321754 348222 324334 354174
rect 321754 346544 322334 348222
rect 323754 346544 324334 348222
rect 321754 345900 324334 346544
rect 411754 355098 414334 355446
rect 411754 354174 412604 355098
rect 413280 354174 414334 355098
rect 411754 348222 414334 354174
rect 411754 346544 412334 348222
rect 413754 346544 414334 348222
rect 411754 345900 414334 346544
rect 501754 355098 504334 355446
rect 501754 354174 502604 355098
rect 503280 354174 504334 355098
rect 501754 348222 504334 354174
rect 501754 346544 502334 348222
rect 503754 346544 504334 348222
rect 501754 345900 504334 346544
rect 63816 276794 66396 277438
rect 63816 275116 64332 276794
rect 65752 275116 66396 276794
rect 63816 269424 66396 275116
rect 63816 268500 64750 269424
rect 65426 268500 66396 269424
rect 63816 267892 66396 268500
rect 152940 276590 155520 277234
rect 152940 274912 153456 276590
rect 154876 274912 155520 276590
rect 152940 269220 155520 274912
rect 152940 268296 153874 269220
rect 154550 268296 155520 269220
rect 152940 267688 155520 268296
rect 244194 276402 246774 277046
rect 244194 274724 244710 276402
rect 246130 274724 246774 276402
rect 244194 269032 246774 274724
rect 244194 268108 245128 269032
rect 245804 268108 246774 269032
rect 244194 267500 246774 268108
rect 333816 276794 336396 277438
rect 333816 275116 334332 276794
rect 335752 275116 336396 276794
rect 333816 269424 336396 275116
rect 333816 268500 334750 269424
rect 335426 268500 336396 269424
rect 333816 267892 336396 268500
rect 423816 276794 426396 277438
rect 423816 275116 424332 276794
rect 425752 275116 426396 276794
rect 423816 269424 426396 275116
rect 423816 268500 424750 269424
rect 425426 268500 426396 269424
rect 423816 267892 426396 268500
rect 513816 276794 516396 277438
rect 513816 275116 514332 276794
rect 515752 275116 516396 276794
rect 513816 269424 516396 275116
rect 513816 268500 514750 269424
rect 515426 268500 516396 269424
rect 513816 267892 516396 268500
rect 57138 264800 58098 265040
rect 57138 264320 57258 264800
rect 57978 264320 58098 264800
rect 57138 261380 58098 264320
rect 57138 260600 57318 261380
rect 57978 260600 58098 261380
rect 57138 260240 58098 260600
rect 60858 264800 61818 265040
rect 60858 264320 60978 264800
rect 61698 264320 61818 264800
rect 60858 261380 61818 264320
rect 60858 260600 61038 261380
rect 61698 260600 61818 261380
rect 60858 260240 61818 260600
rect 146262 264596 147222 264836
rect 146262 264116 146382 264596
rect 147102 264116 147222 264596
rect 146262 261176 147222 264116
rect 146262 260396 146442 261176
rect 147102 260396 147222 261176
rect 146262 260036 147222 260396
rect 149982 264596 150942 264836
rect 327138 264800 328098 265040
rect 149982 264116 150102 264596
rect 150822 264116 150942 264596
rect 149982 261176 150942 264116
rect 149982 260396 150162 261176
rect 150822 260396 150942 261176
rect 149982 260036 150942 260396
rect 237516 264408 238476 264648
rect 237516 263928 237636 264408
rect 238356 263928 238476 264408
rect 237516 260988 238476 263928
rect 237516 260208 237696 260988
rect 238356 260208 238476 260988
rect 237516 259848 238476 260208
rect 241236 264408 242196 264648
rect 241236 263928 241356 264408
rect 242076 263928 242196 264408
rect 241236 260988 242196 263928
rect 241236 260208 241416 260988
rect 242076 260208 242196 260988
rect 327138 264320 327258 264800
rect 327978 264320 328098 264800
rect 327138 261380 328098 264320
rect 327138 260600 327318 261380
rect 327978 260600 328098 261380
rect 327138 260240 328098 260600
rect 330858 264800 331818 265040
rect 330858 264320 330978 264800
rect 331698 264320 331818 264800
rect 330858 261380 331818 264320
rect 330858 260600 331038 261380
rect 331698 260600 331818 261380
rect 330858 260240 331818 260600
rect 417138 264800 418098 265040
rect 417138 264320 417258 264800
rect 417978 264320 418098 264800
rect 417138 261380 418098 264320
rect 417138 260600 417318 261380
rect 417978 260600 418098 261380
rect 417138 260240 418098 260600
rect 420858 264800 421818 265040
rect 420858 264320 420978 264800
rect 421698 264320 421818 264800
rect 420858 261380 421818 264320
rect 420858 260600 421038 261380
rect 421698 260600 421818 261380
rect 420858 260240 421818 260600
rect 507138 264800 508098 265040
rect 507138 264320 507258 264800
rect 507978 264320 508098 264800
rect 507138 261380 508098 264320
rect 507138 260600 507318 261380
rect 507978 260600 508098 261380
rect 507138 260240 508098 260600
rect 510858 264800 511818 265040
rect 510858 264320 510978 264800
rect 511698 264320 511818 264800
rect 510858 261380 511818 264320
rect 510858 260600 511038 261380
rect 511698 260600 511818 261380
rect 510858 260240 511818 260600
rect 241236 259848 242196 260208
rect 319050 254443 320000 254444
rect 317669 253495 319051 254443
rect 319999 253495 320000 254443
rect 53160 251360 56122 252058
rect 53160 251040 53194 251360
rect 53514 251300 56122 251360
rect 53514 251100 55884 251300
rect 56084 251100 56122 251300
rect 53514 251040 56122 251100
rect 53160 250732 56122 251040
rect 63742 251955 67282 252040
rect 230652 251962 230980 251963
rect 63742 251824 67291 251955
rect 63742 251540 66566 251824
rect 63742 251090 63948 251540
rect 64398 251190 66566 251540
rect 67218 251190 67291 251824
rect 64398 251090 67291 251190
rect 63742 251079 67291 251090
rect 142284 251156 145246 251854
rect 63742 250770 67282 251079
rect 142284 250836 142318 251156
rect 142638 251096 145246 251156
rect 142638 250896 145008 251096
rect 145208 250896 145246 251096
rect 142638 250836 145246 250896
rect 142284 250528 145246 250836
rect 152866 251751 156406 251836
rect 152866 251620 156415 251751
rect 152866 251336 155690 251620
rect 152866 250886 153072 251336
rect 153522 250986 155690 251336
rect 156342 250986 156415 251620
rect 230005 251636 230653 251962
rect 230979 251636 230980 251962
rect 230005 251357 230331 251636
rect 230652 251635 230980 251636
rect 317669 251774 318617 253495
rect 319050 253494 320000 253495
rect 250746 251308 251170 251309
rect 153522 250886 156415 250986
rect 152866 250875 156415 250886
rect 250746 250886 250747 251308
rect 251169 250886 251783 251308
rect 250746 250885 251170 250886
rect 152866 250566 156406 250875
rect 339825 248090 341326 250662
rect 339824 248089 341327 248090
rect 339824 246588 339825 248089
rect 341326 246588 341327 248089
rect 409662 247805 410754 247806
rect 409662 246715 409663 247805
rect 410753 246715 410754 247805
rect 499662 247805 500754 247806
rect 409662 246714 410754 246715
rect 428317 247410 429189 247411
rect 339824 246587 341327 246588
rect 409663 245900 410753 246714
rect 428317 246540 428318 247410
rect 429188 246540 430183 247410
rect 499662 246715 499663 247805
rect 500753 246715 500754 247805
rect 499662 246714 500754 246715
rect 518317 247410 519189 247411
rect 428317 246539 429189 246540
rect 499663 245900 500753 246714
rect 518317 246540 518318 247410
rect 519188 246540 520183 247410
rect 518317 246539 519189 246540
rect 57078 243020 58038 243380
rect 57078 242240 57258 243020
rect 57918 242240 58038 243020
rect 57078 239300 58038 242240
rect 57078 238820 57198 239300
rect 57918 238820 58038 239300
rect 57078 238580 58038 238820
rect 60798 243020 61758 243380
rect 60798 242240 60978 243020
rect 61638 242240 61758 243020
rect 60798 239300 61758 242240
rect 60798 238820 60918 239300
rect 61638 238820 61758 239300
rect 60798 238580 61758 238820
rect 146202 242816 147162 243176
rect 146202 242036 146382 242816
rect 147042 242036 147162 242816
rect 146202 239096 147162 242036
rect 146202 238616 146322 239096
rect 147042 238616 147162 239096
rect 146202 238376 147162 238616
rect 149922 242816 150882 243176
rect 327078 243020 328038 243380
rect 149922 242036 150102 242816
rect 150762 242036 150882 242816
rect 149922 239096 150882 242036
rect 149922 238616 150042 239096
rect 150762 238616 150882 239096
rect 149922 238376 150882 238616
rect 237456 242628 238416 242988
rect 237456 241848 237636 242628
rect 238296 241848 238416 242628
rect 237456 238908 238416 241848
rect 237456 238428 237576 238908
rect 238296 238428 238416 238908
rect 237456 238188 238416 238428
rect 241176 242628 242136 242988
rect 241176 241848 241356 242628
rect 242016 241848 242136 242628
rect 241176 238908 242136 241848
rect 241176 238428 241296 238908
rect 242016 238428 242136 238908
rect 327078 242240 327258 243020
rect 327918 242240 328038 243020
rect 327078 239300 328038 242240
rect 327078 238820 327198 239300
rect 327918 238820 328038 239300
rect 327078 238580 328038 238820
rect 330798 243020 331758 243380
rect 330798 242240 330978 243020
rect 331638 242240 331758 243020
rect 330798 239300 331758 242240
rect 330798 238820 330918 239300
rect 331638 238820 331758 239300
rect 330798 238580 331758 238820
rect 417078 243020 418038 243380
rect 417078 242240 417258 243020
rect 417918 242240 418038 243020
rect 417078 239300 418038 242240
rect 417078 238820 417198 239300
rect 417918 238820 418038 239300
rect 417078 238580 418038 238820
rect 420798 243020 421758 243380
rect 420798 242240 420978 243020
rect 421638 242240 421758 243020
rect 420798 239300 421758 242240
rect 420798 238820 420918 239300
rect 421638 238820 421758 239300
rect 420798 238580 421758 238820
rect 507078 243020 508038 243380
rect 507078 242240 507258 243020
rect 507918 242240 508038 243020
rect 507078 239300 508038 242240
rect 507078 238820 507198 239300
rect 507918 238820 508038 239300
rect 507078 238580 508038 238820
rect 510798 243020 511758 243380
rect 510798 242240 510978 243020
rect 511638 242240 511758 243020
rect 510798 239300 511758 242240
rect 510798 238820 510918 239300
rect 511638 238820 511758 239300
rect 510798 238580 511758 238820
rect 241176 238188 242136 238428
rect 51754 235098 54334 235446
rect 51754 234174 52604 235098
rect 53280 234174 54334 235098
rect 51754 228222 54334 234174
rect 51754 226544 52334 228222
rect 53754 226544 54334 228222
rect 51754 225900 54334 226544
rect 140878 234894 143458 235242
rect 321754 235098 324334 235446
rect 140878 233970 141728 234894
rect 142404 233970 143458 234894
rect 140878 228018 143458 233970
rect 140878 226340 141458 228018
rect 142878 226340 143458 228018
rect 140878 225696 143458 226340
rect 232132 234706 234712 235054
rect 232132 233782 232982 234706
rect 233658 233782 234712 234706
rect 232132 227830 234712 233782
rect 232132 226152 232712 227830
rect 234132 226152 234712 227830
rect 232132 225508 234712 226152
rect 321754 234174 322604 235098
rect 323280 234174 324334 235098
rect 321754 228222 324334 234174
rect 321754 226544 322334 228222
rect 323754 226544 324334 228222
rect 321754 225900 324334 226544
rect 411754 235098 414334 235446
rect 411754 234174 412604 235098
rect 413280 234174 414334 235098
rect 411754 228222 414334 234174
rect 411754 226544 412334 228222
rect 413754 226544 414334 228222
rect 411754 225900 414334 226544
rect 501754 235098 504334 235446
rect 501754 234174 502604 235098
rect 503280 234174 504334 235098
rect 501754 228222 504334 234174
rect 501754 226544 502334 228222
rect 503754 226544 504334 228222
rect 501754 225900 504334 226544
rect 57138 158700 58098 158940
rect 57138 158220 57258 158700
rect 57978 158220 58098 158700
rect 57138 155280 58098 158220
rect 57138 154500 57318 155280
rect 57978 154500 58098 155280
rect 57138 154140 58098 154500
rect 60858 158700 61818 158940
rect 60858 158220 60978 158700
rect 61698 158220 61818 158700
rect 60858 155280 61818 158220
rect 60858 154500 61038 155280
rect 61698 154500 61818 155280
rect 60858 154140 61818 154500
rect 147138 158700 148098 158940
rect 147138 158220 147258 158700
rect 147978 158220 148098 158700
rect 147138 155280 148098 158220
rect 147138 154500 147318 155280
rect 147978 154500 148098 155280
rect 147138 154140 148098 154500
rect 150858 158700 151818 158940
rect 150858 158220 150978 158700
rect 151698 158220 151818 158700
rect 150858 155280 151818 158220
rect 150858 154500 151038 155280
rect 151698 154500 151818 155280
rect 150858 154140 151818 154500
rect 237138 158700 238098 158940
rect 237138 158220 237258 158700
rect 237978 158220 238098 158700
rect 237138 155280 238098 158220
rect 237138 154500 237318 155280
rect 237978 154500 238098 155280
rect 237138 154140 238098 154500
rect 240858 158700 241818 158940
rect 240858 158220 240978 158700
rect 241698 158220 241818 158700
rect 240858 155280 241818 158220
rect 240858 154500 241038 155280
rect 241698 154500 241818 155280
rect 240858 154140 241818 154500
rect 327138 158700 328098 158940
rect 327138 158220 327258 158700
rect 327978 158220 328098 158700
rect 327138 155280 328098 158220
rect 327138 154500 327318 155280
rect 327978 154500 328098 155280
rect 327138 154140 328098 154500
rect 330858 158700 331818 158940
rect 330858 158220 330978 158700
rect 331698 158220 331818 158700
rect 330858 155280 331818 158220
rect 330858 154500 331038 155280
rect 331698 154500 331818 155280
rect 330858 154140 331818 154500
rect 417138 158700 418098 158940
rect 417138 158220 417258 158700
rect 417978 158220 418098 158700
rect 417138 155280 418098 158220
rect 417138 154500 417318 155280
rect 417978 154500 418098 155280
rect 417138 154140 418098 154500
rect 420858 158700 421818 158940
rect 420858 158220 420978 158700
rect 421698 158220 421818 158700
rect 420858 155280 421818 158220
rect 420858 154500 421038 155280
rect 421698 154500 421818 155280
rect 420858 154140 421818 154500
rect 507138 158700 508098 158940
rect 507138 158220 507258 158700
rect 507978 158220 508098 158700
rect 507138 155280 508098 158220
rect 507138 154500 507318 155280
rect 507978 154500 508098 155280
rect 507138 154140 508098 154500
rect 510858 158700 511818 158940
rect 510858 158220 510978 158700
rect 511698 158220 511818 158700
rect 510858 155280 511818 158220
rect 510858 154500 511038 155280
rect 511698 154500 511818 155280
rect 510858 154140 511818 154500
rect 53160 145260 56122 145958
rect 53160 144940 53194 145260
rect 53514 145200 56122 145260
rect 53514 145000 55884 145200
rect 56084 145000 56122 145200
rect 53514 144940 56122 145000
rect 53160 144632 56122 144940
rect 63742 145855 67282 145940
rect 63742 145724 67291 145855
rect 63742 145440 66566 145724
rect 63742 144990 63948 145440
rect 64398 145090 66566 145440
rect 67218 145090 67291 145724
rect 64398 144990 67291 145090
rect 63742 144979 67291 144990
rect 143160 145260 146122 145958
rect 63742 144670 67282 144979
rect 143160 144940 143194 145260
rect 143514 145200 146122 145260
rect 143514 145000 145884 145200
rect 146084 145000 146122 145200
rect 143514 144940 146122 145000
rect 143160 144632 146122 144940
rect 153742 145855 157282 145940
rect 153742 145724 157291 145855
rect 153742 145440 156566 145724
rect 153742 144990 153948 145440
rect 154398 145090 156566 145440
rect 157218 145090 157291 145724
rect 154398 144990 157291 145090
rect 153742 144979 157291 144990
rect 233160 145260 236122 145958
rect 153742 144670 157282 144979
rect 233160 144940 233194 145260
rect 233514 145200 236122 145260
rect 233514 145000 235884 145200
rect 236084 145000 236122 145200
rect 233514 144940 236122 145000
rect 233160 144632 236122 144940
rect 243742 145855 247282 145940
rect 243742 145724 247291 145855
rect 243742 145440 246566 145724
rect 243742 144990 243948 145440
rect 244398 145090 246566 145440
rect 247218 145090 247291 145724
rect 244398 144990 247291 145090
rect 243742 144979 247291 144990
rect 323160 145260 326122 145958
rect 243742 144670 247282 144979
rect 323160 144940 323194 145260
rect 323514 145200 326122 145260
rect 323514 145000 325884 145200
rect 326084 145000 326122 145200
rect 323514 144940 326122 145000
rect 323160 144632 326122 144940
rect 333742 145855 337282 145940
rect 333742 145724 337291 145855
rect 333742 145440 336566 145724
rect 333742 144990 333948 145440
rect 334398 145090 336566 145440
rect 337218 145090 337291 145724
rect 334398 144990 337291 145090
rect 333742 144979 337291 144990
rect 413160 145260 416122 145958
rect 333742 144670 337282 144979
rect 413160 144940 413194 145260
rect 413514 145200 416122 145260
rect 413514 145000 415884 145200
rect 416084 145000 416122 145200
rect 413514 144940 416122 145000
rect 413160 144632 416122 144940
rect 423742 145855 427282 145940
rect 423742 145724 427291 145855
rect 423742 145440 426566 145724
rect 423742 144990 423948 145440
rect 424398 145090 426566 145440
rect 427218 145090 427291 145724
rect 424398 144990 427291 145090
rect 423742 144979 427291 144990
rect 503160 145260 506122 145958
rect 423742 144670 427282 144979
rect 503160 144940 503194 145260
rect 503514 145200 506122 145260
rect 503514 145000 505884 145200
rect 506084 145000 506122 145200
rect 503514 144940 506122 145000
rect 503160 144632 506122 144940
rect 513742 145855 517282 145940
rect 513742 145724 517291 145855
rect 513742 145440 516566 145724
rect 513742 144990 513948 145440
rect 514398 145090 516566 145440
rect 517218 145090 517291 145724
rect 514398 144990 517291 145090
rect 513742 144979 517291 144990
rect 513742 144670 517282 144979
rect 57078 136920 58038 137280
rect 57078 136140 57258 136920
rect 57918 136140 58038 136920
rect 57078 133200 58038 136140
rect 57078 132720 57198 133200
rect 57918 132720 58038 133200
rect 57078 132480 58038 132720
rect 60798 136920 61758 137280
rect 60798 136140 60978 136920
rect 61638 136140 61758 136920
rect 60798 133200 61758 136140
rect 60798 132720 60918 133200
rect 61638 132720 61758 133200
rect 60798 132480 61758 132720
rect 147078 136920 148038 137280
rect 147078 136140 147258 136920
rect 147918 136140 148038 136920
rect 147078 133200 148038 136140
rect 147078 132720 147198 133200
rect 147918 132720 148038 133200
rect 147078 132480 148038 132720
rect 150798 136920 151758 137280
rect 150798 136140 150978 136920
rect 151638 136140 151758 136920
rect 150798 133200 151758 136140
rect 150798 132720 150918 133200
rect 151638 132720 151758 133200
rect 150798 132480 151758 132720
rect 237078 136920 238038 137280
rect 237078 136140 237258 136920
rect 237918 136140 238038 136920
rect 237078 133200 238038 136140
rect 237078 132720 237198 133200
rect 237918 132720 238038 133200
rect 237078 132480 238038 132720
rect 240798 136920 241758 137280
rect 240798 136140 240978 136920
rect 241638 136140 241758 136920
rect 240798 133200 241758 136140
rect 240798 132720 240918 133200
rect 241638 132720 241758 133200
rect 240798 132480 241758 132720
rect 327078 136920 328038 137280
rect 327078 136140 327258 136920
rect 327918 136140 328038 136920
rect 327078 133200 328038 136140
rect 327078 132720 327198 133200
rect 327918 132720 328038 133200
rect 327078 132480 328038 132720
rect 330798 136920 331758 137280
rect 330798 136140 330978 136920
rect 331638 136140 331758 136920
rect 330798 133200 331758 136140
rect 330798 132720 330918 133200
rect 331638 132720 331758 133200
rect 330798 132480 331758 132720
rect 417078 136920 418038 137280
rect 417078 136140 417258 136920
rect 417918 136140 418038 136920
rect 417078 133200 418038 136140
rect 417078 132720 417198 133200
rect 417918 132720 418038 133200
rect 417078 132480 418038 132720
rect 420798 136920 421758 137280
rect 420798 136140 420978 136920
rect 421638 136140 421758 136920
rect 420798 133200 421758 136140
rect 420798 132720 420918 133200
rect 421638 132720 421758 133200
rect 420798 132480 421758 132720
rect 507078 136920 508038 137280
rect 507078 136140 507258 136920
rect 507918 136140 508038 136920
rect 507078 133200 508038 136140
rect 507078 132720 507198 133200
rect 507918 132720 508038 133200
rect 507078 132480 508038 132720
rect 510798 136920 511758 137280
rect 510798 136140 510978 136920
rect 511638 136140 511758 136920
rect 510798 133200 511758 136140
rect 510798 132720 510918 133200
rect 511638 132720 511758 133200
rect 510798 132480 511758 132720
rect 57138 68700 58098 68940
rect 57138 68220 57258 68700
rect 57978 68220 58098 68700
rect 57138 65280 58098 68220
rect 57138 64500 57318 65280
rect 57978 64500 58098 65280
rect 57138 64140 58098 64500
rect 60858 68700 61818 68940
rect 60858 68220 60978 68700
rect 61698 68220 61818 68700
rect 60858 65280 61818 68220
rect 60858 64500 61038 65280
rect 61698 64500 61818 65280
rect 60858 64140 61818 64500
rect 147138 68700 148098 68940
rect 147138 68220 147258 68700
rect 147978 68220 148098 68700
rect 147138 65280 148098 68220
rect 147138 64500 147318 65280
rect 147978 64500 148098 65280
rect 147138 64140 148098 64500
rect 150858 68700 151818 68940
rect 150858 68220 150978 68700
rect 151698 68220 151818 68700
rect 150858 65280 151818 68220
rect 150858 64500 151038 65280
rect 151698 64500 151818 65280
rect 150858 64140 151818 64500
rect 237138 68700 238098 68940
rect 237138 68220 237258 68700
rect 237978 68220 238098 68700
rect 237138 65280 238098 68220
rect 237138 64500 237318 65280
rect 237978 64500 238098 65280
rect 237138 64140 238098 64500
rect 240858 68700 241818 68940
rect 240858 68220 240978 68700
rect 241698 68220 241818 68700
rect 240858 65280 241818 68220
rect 240858 64500 241038 65280
rect 241698 64500 241818 65280
rect 240858 64140 241818 64500
rect 327138 68700 328098 68940
rect 327138 68220 327258 68700
rect 327978 68220 328098 68700
rect 327138 65280 328098 68220
rect 327138 64500 327318 65280
rect 327978 64500 328098 65280
rect 327138 64140 328098 64500
rect 330858 68700 331818 68940
rect 330858 68220 330978 68700
rect 331698 68220 331818 68700
rect 330858 65280 331818 68220
rect 330858 64500 331038 65280
rect 331698 64500 331818 65280
rect 330858 64140 331818 64500
rect 417138 68700 418098 68940
rect 417138 68220 417258 68700
rect 417978 68220 418098 68700
rect 417138 65280 418098 68220
rect 417138 64500 417318 65280
rect 417978 64500 418098 65280
rect 417138 64140 418098 64500
rect 420858 68700 421818 68940
rect 420858 68220 420978 68700
rect 421698 68220 421818 68700
rect 420858 65280 421818 68220
rect 420858 64500 421038 65280
rect 421698 64500 421818 65280
rect 420858 64140 421818 64500
rect 507138 68700 508098 68940
rect 507138 68220 507258 68700
rect 507978 68220 508098 68700
rect 507138 65280 508098 68220
rect 507138 64500 507318 65280
rect 507978 64500 508098 65280
rect 507138 64140 508098 64500
rect 510858 68700 511818 68940
rect 510858 68220 510978 68700
rect 511698 68220 511818 68700
rect 510858 65280 511818 68220
rect 510858 64500 511038 65280
rect 511698 64500 511818 65280
rect 510858 64140 511818 64500
rect 53160 55260 56122 55958
rect 53160 54940 53194 55260
rect 53514 55200 56122 55260
rect 53514 55000 55884 55200
rect 56084 55000 56122 55200
rect 53514 54940 56122 55000
rect 53160 54632 56122 54940
rect 63742 55855 67282 55940
rect 63742 55724 67291 55855
rect 63742 55440 66566 55724
rect 63742 54990 63948 55440
rect 64398 55090 66566 55440
rect 67218 55090 67291 55724
rect 64398 54990 67291 55090
rect 63742 54979 67291 54990
rect 143160 55260 146122 55958
rect 63742 54670 67282 54979
rect 143160 54940 143194 55260
rect 143514 55200 146122 55260
rect 143514 55000 145884 55200
rect 146084 55000 146122 55200
rect 143514 54940 146122 55000
rect 143160 54632 146122 54940
rect 153742 55855 157282 55940
rect 153742 55724 157291 55855
rect 153742 55440 156566 55724
rect 153742 54990 153948 55440
rect 154398 55090 156566 55440
rect 157218 55090 157291 55724
rect 154398 54990 157291 55090
rect 153742 54979 157291 54990
rect 233160 55260 236122 55958
rect 153742 54670 157282 54979
rect 233160 54940 233194 55260
rect 233514 55200 236122 55260
rect 233514 55000 235884 55200
rect 236084 55000 236122 55200
rect 233514 54940 236122 55000
rect 233160 54632 236122 54940
rect 243742 55855 247282 55940
rect 243742 55724 247291 55855
rect 243742 55440 246566 55724
rect 243742 54990 243948 55440
rect 244398 55090 246566 55440
rect 247218 55090 247291 55724
rect 244398 54990 247291 55090
rect 243742 54979 247291 54990
rect 323160 55260 326122 55958
rect 243742 54670 247282 54979
rect 323160 54940 323194 55260
rect 323514 55200 326122 55260
rect 323514 55000 325884 55200
rect 326084 55000 326122 55200
rect 323514 54940 326122 55000
rect 323160 54632 326122 54940
rect 333742 55855 337282 55940
rect 333742 55724 337291 55855
rect 333742 55440 336566 55724
rect 333742 54990 333948 55440
rect 334398 55090 336566 55440
rect 337218 55090 337291 55724
rect 334398 54990 337291 55090
rect 333742 54979 337291 54990
rect 413160 55260 416122 55958
rect 333742 54670 337282 54979
rect 413160 54940 413194 55260
rect 413514 55200 416122 55260
rect 413514 55000 415884 55200
rect 416084 55000 416122 55200
rect 413514 54940 416122 55000
rect 413160 54632 416122 54940
rect 423742 55855 427282 55940
rect 423742 55724 427291 55855
rect 423742 55440 426566 55724
rect 423742 54990 423948 55440
rect 424398 55090 426566 55440
rect 427218 55090 427291 55724
rect 424398 54990 427291 55090
rect 423742 54979 427291 54990
rect 503160 55260 506122 55958
rect 423742 54670 427282 54979
rect 503160 54940 503194 55260
rect 503514 55200 506122 55260
rect 503514 55000 505884 55200
rect 506084 55000 506122 55200
rect 503514 54940 506122 55000
rect 503160 54632 506122 54940
rect 513742 55855 517282 55940
rect 513742 55724 517291 55855
rect 513742 55440 516566 55724
rect 513742 54990 513948 55440
rect 514398 55090 516566 55440
rect 517218 55090 517291 55724
rect 514398 54990 517291 55090
rect 513742 54979 517291 54990
rect 513742 54670 517282 54979
rect 57078 46920 58038 47280
rect 57078 46140 57258 46920
rect 57918 46140 58038 46920
rect 57078 43200 58038 46140
rect 57078 42720 57198 43200
rect 57918 42720 58038 43200
rect 57078 42480 58038 42720
rect 60798 46920 61758 47280
rect 60798 46140 60978 46920
rect 61638 46140 61758 46920
rect 60798 43200 61758 46140
rect 60798 42720 60918 43200
rect 61638 42720 61758 43200
rect 60798 42480 61758 42720
rect 147078 46920 148038 47280
rect 147078 46140 147258 46920
rect 147918 46140 148038 46920
rect 147078 43200 148038 46140
rect 147078 42720 147198 43200
rect 147918 42720 148038 43200
rect 147078 42480 148038 42720
rect 150798 46920 151758 47280
rect 150798 46140 150978 46920
rect 151638 46140 151758 46920
rect 150798 43200 151758 46140
rect 150798 42720 150918 43200
rect 151638 42720 151758 43200
rect 150798 42480 151758 42720
rect 237078 46920 238038 47280
rect 237078 46140 237258 46920
rect 237918 46140 238038 46920
rect 237078 43200 238038 46140
rect 237078 42720 237198 43200
rect 237918 42720 238038 43200
rect 237078 42480 238038 42720
rect 240798 46920 241758 47280
rect 240798 46140 240978 46920
rect 241638 46140 241758 46920
rect 240798 43200 241758 46140
rect 240798 42720 240918 43200
rect 241638 42720 241758 43200
rect 240798 42480 241758 42720
rect 327078 46920 328038 47280
rect 327078 46140 327258 46920
rect 327918 46140 328038 46920
rect 327078 43200 328038 46140
rect 327078 42720 327198 43200
rect 327918 42720 328038 43200
rect 327078 42480 328038 42720
rect 330798 46920 331758 47280
rect 330798 46140 330978 46920
rect 331638 46140 331758 46920
rect 330798 43200 331758 46140
rect 330798 42720 330918 43200
rect 331638 42720 331758 43200
rect 330798 42480 331758 42720
rect 417078 46920 418038 47280
rect 417078 46140 417258 46920
rect 417918 46140 418038 46920
rect 417078 43200 418038 46140
rect 417078 42720 417198 43200
rect 417918 42720 418038 43200
rect 417078 42480 418038 42720
rect 420798 46920 421758 47280
rect 420798 46140 420978 46920
rect 421638 46140 421758 46920
rect 420798 43200 421758 46140
rect 420798 42720 420918 43200
rect 421638 42720 421758 43200
rect 420798 42480 421758 42720
rect 507078 46920 508038 47280
rect 507078 46140 507258 46920
rect 507918 46140 508038 46920
rect 507078 43200 508038 46140
rect 507078 42720 507198 43200
rect 507918 42720 508038 43200
rect 507078 42480 508038 42720
rect 510798 46920 511758 47280
rect 510798 46140 510978 46920
rect 511638 46140 511758 46920
rect 510798 43200 511758 46140
rect 510798 42720 510918 43200
rect 511638 42720 511758 43200
rect 510798 42480 511758 42720
<< via4 >>
rect 327060 670144 327780 670624
rect 57258 668220 57978 668700
rect 60978 668220 61698 668700
rect 147258 668220 147978 668700
rect 150978 668220 151698 668700
rect 237258 668220 237978 668700
rect 240978 668220 241698 668700
rect 330780 670144 331500 670624
rect 417060 670144 417780 670624
rect 420780 670144 421500 670624
rect 507060 670144 507780 670624
rect 510780 670144 511500 670624
rect 322996 656864 323316 657184
rect 336368 657014 337020 657648
rect 412996 656864 413316 657184
rect 426368 657014 427020 657648
rect 502996 656864 503316 657184
rect 516368 657014 517020 657648
rect 53194 654940 53514 655260
rect 66566 655090 67218 655724
rect 143194 654940 143514 655260
rect 156566 655090 157218 655724
rect 233194 654940 233514 655260
rect 246566 655090 247218 655724
rect 57198 642720 57918 643200
rect 60918 642720 61638 643200
rect 147198 642720 147918 643200
rect 150918 642720 151638 643200
rect 237198 642720 237918 643200
rect 327000 644644 327720 645124
rect 330720 644644 331440 645124
rect 417000 644644 417720 645124
rect 420720 644644 421440 645124
rect 507000 644644 507720 645124
rect 510720 644644 511440 645124
rect 240918 642720 241638 643200
rect 417060 595144 417780 595624
rect 57258 593220 57978 593700
rect 60978 593220 61698 593700
rect 147258 593220 147978 593700
rect 150978 593220 151698 593700
rect 237258 593220 237978 593700
rect 240978 593220 241698 593700
rect 327258 593220 327978 593700
rect 330978 593220 331698 593700
rect 420780 595144 421500 595624
rect 507060 595144 507780 595624
rect 510780 595144 511500 595624
rect 412996 581864 413316 582184
rect 426368 582014 427020 582648
rect 502996 581864 503316 582184
rect 516368 582014 517020 582648
rect 53194 579940 53514 580260
rect 66566 580090 67218 580724
rect 143194 579940 143514 580260
rect 156566 580090 157218 580724
rect 233194 579940 233514 580260
rect 246566 580090 247218 580724
rect 323194 579940 323514 580260
rect 336566 580090 337218 580724
rect 57198 567720 57918 568200
rect 60918 567720 61638 568200
rect 147198 567720 147918 568200
rect 150918 567720 151638 568200
rect 237198 567720 237918 568200
rect 240918 567720 241638 568200
rect 327198 567720 327918 568200
rect 417000 569644 417720 570124
rect 420720 569644 421440 570124
rect 507000 569644 507720 570124
rect 510720 569644 511440 570124
rect 330918 567720 331638 568200
rect 64332 515116 65752 516794
rect 154332 515116 155752 516794
rect 244332 515116 245752 516794
rect 334332 515116 335752 516794
rect 424332 515116 425752 516794
rect 514332 515116 515752 516794
rect 57258 504320 57978 504800
rect 60978 504320 61698 504800
rect 147258 504320 147978 504800
rect 150978 504320 151698 504800
rect 237258 504320 237978 504800
rect 240978 504320 241698 504800
rect 327258 504320 327978 504800
rect 330978 504320 331698 504800
rect 417258 504320 417978 504800
rect 420978 504320 421698 504800
rect 507258 504320 507978 504800
rect 510978 504320 511698 504800
rect 53194 491040 53514 491360
rect 66566 491190 67218 491824
rect 227669 490826 228617 491774
rect 249825 490662 251326 492163
rect 319627 491423 319953 491749
rect 341405 491278 341827 491700
rect 413194 491040 413514 491360
rect 426566 491190 427218 491824
rect 503194 491040 503514 491360
rect 516566 491190 517218 491824
rect 160183 486540 161053 487410
rect 139663 484810 140753 485900
rect 57198 478820 57918 479300
rect 60918 478820 61638 479300
rect 147198 478820 147918 479300
rect 150918 478820 151638 479300
rect 237198 478820 237918 479300
rect 240918 478820 241638 479300
rect 327198 478820 327918 479300
rect 330918 478820 331638 479300
rect 417198 478820 417918 479300
rect 420918 478820 421638 479300
rect 507198 478820 507918 479300
rect 510918 478820 511638 479300
rect 52334 466544 53754 468222
rect 142334 466544 143754 468222
rect 232334 466544 233754 468222
rect 322334 466544 323754 468222
rect 412334 466544 413754 468222
rect 502334 466544 503754 468222
rect 64332 395116 65752 396794
rect 154332 395116 155752 396794
rect 244332 395116 245752 396794
rect 334332 395116 335752 396794
rect 424332 395116 425752 396794
rect 514332 395116 515752 396794
rect 57258 384320 57978 384800
rect 60978 384320 61698 384800
rect 147258 384320 147978 384800
rect 150978 384320 151698 384800
rect 237258 384320 237978 384800
rect 240978 384320 241698 384800
rect 327258 384320 327978 384800
rect 330978 384320 331698 384800
rect 417258 384320 417978 384800
rect 420978 384320 421698 384800
rect 507258 384320 507978 384800
rect 510978 384320 511698 384800
rect 227669 370826 228617 371774
rect 249825 370662 251326 372163
rect 319627 371423 319953 371749
rect 341405 371278 341827 371700
rect 413194 371040 413514 371360
rect 426566 371190 427218 371824
rect 503194 371040 503514 371360
rect 516566 371190 517218 371824
rect 70183 366540 71053 367410
rect 49663 364810 50753 365900
rect 160183 366540 161053 367410
rect 139663 364810 140753 365900
rect 57198 358820 57918 359300
rect 60918 358820 61638 359300
rect 147198 358820 147918 359300
rect 150918 358820 151638 359300
rect 237198 358820 237918 359300
rect 240918 358820 241638 359300
rect 327198 358820 327918 359300
rect 330918 358820 331638 359300
rect 417198 358820 417918 359300
rect 420918 358820 421638 359300
rect 507198 358820 507918 359300
rect 510918 358820 511638 359300
rect 52334 346544 53754 348222
rect 142334 346544 143754 348222
rect 232334 346544 233754 348222
rect 322334 346544 323754 348222
rect 412334 346544 413754 348222
rect 502334 346544 503754 348222
rect 64332 275116 65752 276794
rect 153456 274912 154876 276590
rect 244710 274724 246130 276402
rect 334332 275116 335752 276794
rect 424332 275116 425752 276794
rect 514332 275116 515752 276794
rect 57258 264320 57978 264800
rect 60978 264320 61698 264800
rect 146382 264116 147102 264596
rect 150102 264116 150822 264596
rect 237636 263928 238356 264408
rect 241356 263928 242076 264408
rect 327258 264320 327978 264800
rect 330978 264320 331698 264800
rect 417258 264320 417978 264800
rect 420978 264320 421698 264800
rect 507258 264320 507978 264800
rect 510978 264320 511698 264800
rect 53194 251040 53514 251360
rect 66566 251190 67218 251824
rect 142318 250836 142638 251156
rect 155690 250986 156342 251620
rect 230005 251031 230331 251357
rect 251783 250886 252205 251308
rect 317669 250826 318617 251774
rect 339825 250662 341326 252163
rect 430183 246540 431053 247410
rect 409663 244810 410753 245900
rect 520183 246540 521053 247410
rect 499663 244810 500753 245900
rect 57198 238820 57918 239300
rect 60918 238820 61638 239300
rect 146322 238616 147042 239096
rect 150042 238616 150762 239096
rect 237576 238428 238296 238908
rect 241296 238428 242016 238908
rect 327198 238820 327918 239300
rect 330918 238820 331638 239300
rect 417198 238820 417918 239300
rect 420918 238820 421638 239300
rect 507198 238820 507918 239300
rect 510918 238820 511638 239300
rect 52334 226544 53754 228222
rect 141458 226340 142878 228018
rect 232712 226152 234132 227830
rect 322334 226544 323754 228222
rect 412334 226544 413754 228222
rect 502334 226544 503754 228222
rect 57258 158220 57978 158700
rect 60978 158220 61698 158700
rect 147258 158220 147978 158700
rect 150978 158220 151698 158700
rect 237258 158220 237978 158700
rect 240978 158220 241698 158700
rect 327258 158220 327978 158700
rect 330978 158220 331698 158700
rect 417258 158220 417978 158700
rect 420978 158220 421698 158700
rect 507258 158220 507978 158700
rect 510978 158220 511698 158700
rect 53194 144940 53514 145260
rect 66566 145090 67218 145724
rect 143194 144940 143514 145260
rect 156566 145090 157218 145724
rect 233194 144940 233514 145260
rect 246566 145090 247218 145724
rect 323194 144940 323514 145260
rect 336566 145090 337218 145724
rect 413194 144940 413514 145260
rect 426566 145090 427218 145724
rect 503194 144940 503514 145260
rect 516566 145090 517218 145724
rect 57198 132720 57918 133200
rect 60918 132720 61638 133200
rect 147198 132720 147918 133200
rect 150918 132720 151638 133200
rect 237198 132720 237918 133200
rect 240918 132720 241638 133200
rect 327198 132720 327918 133200
rect 330918 132720 331638 133200
rect 417198 132720 417918 133200
rect 420918 132720 421638 133200
rect 507198 132720 507918 133200
rect 510918 132720 511638 133200
rect 57258 68220 57978 68700
rect 60978 68220 61698 68700
rect 147258 68220 147978 68700
rect 150978 68220 151698 68700
rect 237258 68220 237978 68700
rect 240978 68220 241698 68700
rect 327258 68220 327978 68700
rect 330978 68220 331698 68700
rect 417258 68220 417978 68700
rect 420978 68220 421698 68700
rect 507258 68220 507978 68700
rect 510978 68220 511698 68700
rect 53194 54940 53514 55260
rect 66566 55090 67218 55724
rect 143194 54940 143514 55260
rect 156566 55090 157218 55724
rect 233194 54940 233514 55260
rect 246566 55090 247218 55724
rect 323194 54940 323514 55260
rect 336566 55090 337218 55724
rect 413194 54940 413514 55260
rect 426566 55090 427218 55724
rect 503194 54940 503514 55260
rect 516566 55090 517218 55724
rect 57198 42720 57918 43200
rect 60918 42720 61638 43200
rect 147198 42720 147918 43200
rect 150918 42720 151638 43200
rect 237198 42720 237918 43200
rect 240918 42720 241638 43200
rect 327198 42720 327918 43200
rect 330918 42720 331638 43200
rect 417198 42720 417918 43200
rect 420918 42720 421638 43200
rect 507198 42720 507918 43200
rect 510918 42720 511638 43200
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 30332 676200 46332 681820
rect 30332 674940 58098 676200
rect 73518 676140 89518 681840
rect 72558 676124 89518 676140
rect 60790 675008 89518 676124
rect 60790 674992 63836 675008
rect 72558 675000 89518 675008
rect 30332 673040 46332 674940
rect 30198 672040 46338 673040
rect 30332 665620 46332 672040
rect 57124 669120 58092 674940
rect 57104 668700 58114 669120
rect 57104 668220 57258 668700
rect 57978 668220 58114 668700
rect 57104 668020 58114 668220
rect 60824 668700 61834 674992
rect 60824 668220 60978 668700
rect 61698 668220 61834 668700
rect 60824 668020 61834 668220
rect 73518 665640 89518 675000
rect 120332 676200 136332 681820
rect 120332 674940 148098 676200
rect 163518 676140 179518 681840
rect 162558 676124 179518 676140
rect 150790 675008 179518 676124
rect 150790 674992 153836 675008
rect 162558 675000 179518 675008
rect 120332 673040 136332 674940
rect 120198 672040 136338 673040
rect 120332 665620 136332 672040
rect 147124 669120 148092 674940
rect 147104 668700 148114 669120
rect 147104 668220 147258 668700
rect 147978 668220 148114 668700
rect 147104 668020 148114 668220
rect 150824 668700 151834 674992
rect 150824 668220 150978 668700
rect 151698 668220 151834 668700
rect 150824 668020 151834 668220
rect 163518 665640 179518 675000
rect 210332 676200 226332 681820
rect 210332 674940 238098 676200
rect 253518 676140 269518 681840
rect 252558 676124 269518 676140
rect 240790 675008 269518 676124
rect 240790 674992 243836 675008
rect 252558 675000 269518 675008
rect 210332 673040 226332 674940
rect 210198 672040 226338 673040
rect 210332 665620 226332 672040
rect 237124 669120 238092 674940
rect 237104 668700 238114 669120
rect 237104 668220 237258 668700
rect 237978 668220 238114 668700
rect 237104 668020 238114 668220
rect 240824 668700 241834 674992
rect 240824 668220 240978 668700
rect 241698 668220 241834 668700
rect 240824 668020 241834 668220
rect 253518 665640 269518 675000
rect 300134 678124 316134 683744
rect 300134 676864 327900 678124
rect 343320 678064 359320 683764
rect 342360 678048 359320 678064
rect 330592 676932 359320 678048
rect 330592 676916 333638 676932
rect 342360 676924 359320 676932
rect 300134 674964 316134 676864
rect 300000 673964 316140 674964
rect 300134 667544 316134 673964
rect 326926 671044 327894 676864
rect 326906 670624 327916 671044
rect 326906 670144 327060 670624
rect 327780 670144 327916 670624
rect 326906 669944 327916 670144
rect 330626 670624 331636 676916
rect 330626 670144 330780 670624
rect 331500 670144 331636 670624
rect 330626 669944 331636 670144
rect 343320 667564 359320 676924
rect 390134 678124 406134 683744
rect 390134 676864 417900 678124
rect 433320 678064 449320 683764
rect 432360 678048 449320 678064
rect 420592 676932 449320 678048
rect 420592 676916 423638 676932
rect 432360 676924 449320 676932
rect 390134 674964 406134 676864
rect 390000 673964 406140 674964
rect 390134 667544 406134 673964
rect 416926 671044 417894 676864
rect 416906 670624 417916 671044
rect 416906 670144 417060 670624
rect 417780 670144 417916 670624
rect 416906 669944 417916 670144
rect 420626 670624 421636 676916
rect 420626 670144 420780 670624
rect 421500 670144 421636 670624
rect 420626 669944 421636 670144
rect 433320 667564 449320 676924
rect 480134 678124 496134 683744
rect 480134 676864 507900 678124
rect 523320 678064 539320 683764
rect 522360 678048 539320 678064
rect 510592 676932 539320 678048
rect 510592 676916 513638 676932
rect 522360 676924 539320 676932
rect 480134 674964 496134 676864
rect 480000 673964 496140 674964
rect 480134 667544 496134 673964
rect 506926 671044 507894 676864
rect 506906 670624 507916 671044
rect 506906 670144 507060 670624
rect 507780 670144 507916 670624
rect 506906 669944 507916 670144
rect 510626 670624 511636 676916
rect 510626 670144 510780 670624
rect 511500 670144 511636 670624
rect 510626 669944 511636 670144
rect 523320 667564 539320 676924
rect 30398 655954 46398 663140
rect 73428 656094 89428 663106
rect 30398 655950 53488 655954
rect 30398 655260 53546 655950
rect 30398 654940 53194 655260
rect 53514 654940 53546 655260
rect 30398 654664 53546 654940
rect 66398 655724 89428 656094
rect 66398 655090 66566 655724
rect 67218 655090 89428 655724
rect 30398 646940 46398 654664
rect 66398 654554 89428 655090
rect 73428 646906 89428 654554
rect 120398 655954 136398 663140
rect 163428 656094 179428 663106
rect 120398 655950 143488 655954
rect 120398 655260 143546 655950
rect 120398 654940 143194 655260
rect 143514 654940 143546 655260
rect 120398 654664 143546 654940
rect 156398 655724 179428 656094
rect 156398 655090 156566 655724
rect 157218 655090 179428 655724
rect 120398 646940 136398 654664
rect 156398 654554 179428 655090
rect 163428 646906 179428 654554
rect 210398 655954 226398 663140
rect 253428 656094 269428 663106
rect 210398 655950 233488 655954
rect 210398 655260 233546 655950
rect 210398 654940 233194 655260
rect 233514 654940 233546 655260
rect 210398 654664 233546 654940
rect 246398 655724 269428 656094
rect 246398 655090 246566 655724
rect 247218 655090 269428 655724
rect 210398 646940 226398 654664
rect 246398 654554 269428 655090
rect 253428 646906 269428 654554
rect 300200 657878 316200 665064
rect 343230 658018 359230 665030
rect 300200 657874 323290 657878
rect 300200 657184 323348 657874
rect 300200 656864 322996 657184
rect 323316 656864 323348 657184
rect 300200 656588 323348 656864
rect 336200 657648 359230 658018
rect 336200 657014 336368 657648
rect 337020 657014 359230 657648
rect 300200 648864 316200 656588
rect 336200 656478 359230 657014
rect 343230 648830 359230 656478
rect 390200 657878 406200 665064
rect 433230 658018 449230 665030
rect 390200 657874 413290 657878
rect 390200 657184 413348 657874
rect 390200 656864 412996 657184
rect 413316 656864 413348 657184
rect 390200 656588 413348 656864
rect 426200 657648 449230 658018
rect 426200 657014 426368 657648
rect 427020 657014 449230 657648
rect 390200 648864 406200 656588
rect 426200 656478 449230 657014
rect 433230 648830 449230 656478
rect 480200 657878 496200 665064
rect 523230 658018 539230 665030
rect 480200 657874 503290 657878
rect 480200 657184 503348 657874
rect 480200 656864 502996 657184
rect 503316 656864 503348 657184
rect 480200 656588 503348 656864
rect 516200 657648 539230 658018
rect 516200 657014 516368 657648
rect 517020 657014 539230 657648
rect 480200 648864 496200 656588
rect 516200 656478 539230 657014
rect 523230 648830 539230 656478
rect 30318 636264 46318 644418
rect 57044 643200 58054 643400
rect 57044 642720 57198 643200
rect 57918 642720 58054 643200
rect 57044 642300 58054 642720
rect 60764 643200 61774 643400
rect 60764 642720 60918 643200
rect 61638 642720 61774 643200
rect 57064 636264 58032 642300
rect 60764 636428 61774 642720
rect 60730 636412 63776 636428
rect 73428 636412 89428 644276
rect 30318 635338 58072 636264
rect 30318 628218 46318 635338
rect 60730 635296 89428 636412
rect 73400 635188 89428 635296
rect 73428 628076 89428 635188
rect 120318 636264 136318 644418
rect 147044 643200 148054 643400
rect 147044 642720 147198 643200
rect 147918 642720 148054 643200
rect 147044 642300 148054 642720
rect 150764 643200 151774 643400
rect 150764 642720 150918 643200
rect 151638 642720 151774 643200
rect 147064 636264 148032 642300
rect 150764 636428 151774 642720
rect 150730 636412 153776 636428
rect 163428 636412 179428 644276
rect 120318 635338 148072 636264
rect 120318 628218 136318 635338
rect 150730 635296 179428 636412
rect 163400 635188 179428 635296
rect 163428 628076 179428 635188
rect 210318 636264 226318 644418
rect 237044 643200 238054 643400
rect 237044 642720 237198 643200
rect 237918 642720 238054 643200
rect 237044 642300 238054 642720
rect 240764 643200 241774 643400
rect 240764 642720 240918 643200
rect 241638 642720 241774 643200
rect 237064 636264 238032 642300
rect 240764 636428 241774 642720
rect 240730 636412 243776 636428
rect 253428 636412 269428 644276
rect 210318 635338 238072 636264
rect 210318 628218 226318 635338
rect 240730 635296 269428 636412
rect 253400 635188 269428 635296
rect 253428 628076 269428 635188
rect 300120 638188 316120 646342
rect 326846 645124 327856 645324
rect 326846 644644 327000 645124
rect 327720 644644 327856 645124
rect 326846 644224 327856 644644
rect 330566 645124 331576 645324
rect 330566 644644 330720 645124
rect 331440 644644 331576 645124
rect 326866 638188 327834 644224
rect 330566 638352 331576 644644
rect 330532 638336 333578 638352
rect 343230 638336 359230 646200
rect 300120 637262 327874 638188
rect 300120 630142 316120 637262
rect 330532 637220 359230 638336
rect 343202 637112 359230 637220
rect 343230 630000 359230 637112
rect 390120 638188 406120 646342
rect 416846 645124 417856 645324
rect 416846 644644 417000 645124
rect 417720 644644 417856 645124
rect 416846 644224 417856 644644
rect 420566 645124 421576 645324
rect 420566 644644 420720 645124
rect 421440 644644 421576 645124
rect 416866 638188 417834 644224
rect 420566 638352 421576 644644
rect 420532 638336 423578 638352
rect 433230 638336 449230 646200
rect 390120 637262 417874 638188
rect 390120 630142 406120 637262
rect 420532 637220 449230 638336
rect 433202 637112 449230 637220
rect 433230 630000 449230 637112
rect 480120 638188 496120 646342
rect 506846 645124 507856 645324
rect 506846 644644 507000 645124
rect 507720 644644 507856 645124
rect 506846 644224 507856 644644
rect 510566 645124 511576 645324
rect 510566 644644 510720 645124
rect 511440 644644 511576 645124
rect 506866 638188 507834 644224
rect 510566 638352 511576 644644
rect 510532 638336 513578 638352
rect 523230 638336 539230 646200
rect 480120 637262 507874 638188
rect 480120 630142 496120 637262
rect 510532 637220 539230 638336
rect 523202 637112 539230 637220
rect 523230 630000 539230 637112
rect 30332 601200 46332 606820
rect 30332 599940 58098 601200
rect 73518 601140 89518 606840
rect 72558 601124 89518 601140
rect 60790 600008 89518 601124
rect 60790 599992 63836 600008
rect 72558 600000 89518 600008
rect 30332 598040 46332 599940
rect 30198 597040 46338 598040
rect 30332 590620 46332 597040
rect 57124 594120 58092 599940
rect 57104 593700 58114 594120
rect 57104 593220 57258 593700
rect 57978 593220 58114 593700
rect 57104 593020 58114 593220
rect 60824 593700 61834 599992
rect 60824 593220 60978 593700
rect 61698 593220 61834 593700
rect 60824 593020 61834 593220
rect 73518 590640 89518 600000
rect 120332 601200 136332 606820
rect 120332 599940 148098 601200
rect 163518 601140 179518 606840
rect 162558 601124 179518 601140
rect 150790 600008 179518 601124
rect 150790 599992 153836 600008
rect 162558 600000 179518 600008
rect 120332 598040 136332 599940
rect 120198 597040 136338 598040
rect 120332 590620 136332 597040
rect 147124 594120 148092 599940
rect 147104 593700 148114 594120
rect 147104 593220 147258 593700
rect 147978 593220 148114 593700
rect 147104 593020 148114 593220
rect 150824 593700 151834 599992
rect 150824 593220 150978 593700
rect 151698 593220 151834 593700
rect 150824 593020 151834 593220
rect 163518 590640 179518 600000
rect 210332 601200 226332 606820
rect 210332 599940 238098 601200
rect 253518 601140 269518 606840
rect 252558 601124 269518 601140
rect 240790 600008 269518 601124
rect 240790 599992 243836 600008
rect 252558 600000 269518 600008
rect 210332 598040 226332 599940
rect 210198 597040 226338 598040
rect 210332 590620 226332 597040
rect 237124 594120 238092 599940
rect 237104 593700 238114 594120
rect 237104 593220 237258 593700
rect 237978 593220 238114 593700
rect 237104 593020 238114 593220
rect 240824 593700 241834 599992
rect 240824 593220 240978 593700
rect 241698 593220 241834 593700
rect 240824 593020 241834 593220
rect 253518 590640 269518 600000
rect 300332 601200 316332 606820
rect 300332 599940 328098 601200
rect 343518 601140 359518 606840
rect 342558 601124 359518 601140
rect 330790 600008 359518 601124
rect 330790 599992 333836 600008
rect 342558 600000 359518 600008
rect 300332 598040 316332 599940
rect 300198 597040 316338 598040
rect 300332 590620 316332 597040
rect 327124 594120 328092 599940
rect 327104 593700 328114 594120
rect 327104 593220 327258 593700
rect 327978 593220 328114 593700
rect 327104 593020 328114 593220
rect 330824 593700 331834 599992
rect 330824 593220 330978 593700
rect 331698 593220 331834 593700
rect 330824 593020 331834 593220
rect 343518 590640 359518 600000
rect 390134 603124 406134 608744
rect 390134 601864 417900 603124
rect 433320 603064 449320 608764
rect 432360 603048 449320 603064
rect 420592 601932 449320 603048
rect 420592 601916 423638 601932
rect 432360 601924 449320 601932
rect 390134 599964 406134 601864
rect 390000 598964 406140 599964
rect 390134 592544 406134 598964
rect 416926 596044 417894 601864
rect 416906 595624 417916 596044
rect 416906 595144 417060 595624
rect 417780 595144 417916 595624
rect 416906 594944 417916 595144
rect 420626 595624 421636 601916
rect 420626 595144 420780 595624
rect 421500 595144 421636 595624
rect 420626 594944 421636 595144
rect 433320 592564 449320 601924
rect 480134 603124 496134 608744
rect 480134 601864 507900 603124
rect 523320 603064 539320 608764
rect 522360 603048 539320 603064
rect 510592 601932 539320 603048
rect 510592 601916 513638 601932
rect 522360 601924 539320 601932
rect 480134 599964 496134 601864
rect 480000 598964 496140 599964
rect 480134 592544 496134 598964
rect 506926 596044 507894 601864
rect 506906 595624 507916 596044
rect 506906 595144 507060 595624
rect 507780 595144 507916 595624
rect 506906 594944 507916 595144
rect 510626 595624 511636 601916
rect 510626 595144 510780 595624
rect 511500 595144 511636 595624
rect 510626 594944 511636 595144
rect 523320 592564 539320 601924
rect 30398 580954 46398 588140
rect 73428 581094 89428 588106
rect 30398 580950 53488 580954
rect 30398 580260 53546 580950
rect 30398 579940 53194 580260
rect 53514 579940 53546 580260
rect 30398 579664 53546 579940
rect 66398 580724 89428 581094
rect 66398 580090 66566 580724
rect 67218 580090 89428 580724
rect 30398 571940 46398 579664
rect 66398 579554 89428 580090
rect 73428 571906 89428 579554
rect 120398 580954 136398 588140
rect 163428 581094 179428 588106
rect 120398 580950 143488 580954
rect 120398 580260 143546 580950
rect 120398 579940 143194 580260
rect 143514 579940 143546 580260
rect 120398 579664 143546 579940
rect 156398 580724 179428 581094
rect 156398 580090 156566 580724
rect 157218 580090 179428 580724
rect 120398 571940 136398 579664
rect 156398 579554 179428 580090
rect 163428 571906 179428 579554
rect 210398 580954 226398 588140
rect 253428 581094 269428 588106
rect 210398 580950 233488 580954
rect 210398 580260 233546 580950
rect 210398 579940 233194 580260
rect 233514 579940 233546 580260
rect 210398 579664 233546 579940
rect 246398 580724 269428 581094
rect 246398 580090 246566 580724
rect 247218 580090 269428 580724
rect 210398 571940 226398 579664
rect 246398 579554 269428 580090
rect 253428 571906 269428 579554
rect 300398 580954 316398 588140
rect 343428 581094 359428 588106
rect 300398 580950 323488 580954
rect 300398 580260 323546 580950
rect 300398 579940 323194 580260
rect 323514 579940 323546 580260
rect 300398 579664 323546 579940
rect 336398 580724 359428 581094
rect 336398 580090 336566 580724
rect 337218 580090 359428 580724
rect 300398 571940 316398 579664
rect 336398 579554 359428 580090
rect 343428 571906 359428 579554
rect 390200 582878 406200 590064
rect 433230 583018 449230 590030
rect 390200 582874 413290 582878
rect 390200 582184 413348 582874
rect 390200 581864 412996 582184
rect 413316 581864 413348 582184
rect 390200 581588 413348 581864
rect 426200 582648 449230 583018
rect 426200 582014 426368 582648
rect 427020 582014 449230 582648
rect 390200 573864 406200 581588
rect 426200 581478 449230 582014
rect 433230 573830 449230 581478
rect 480200 582878 496200 590064
rect 523230 583018 539230 590030
rect 480200 582874 503290 582878
rect 480200 582184 503348 582874
rect 480200 581864 502996 582184
rect 503316 581864 503348 582184
rect 480200 581588 503348 581864
rect 516200 582648 539230 583018
rect 516200 582014 516368 582648
rect 517020 582014 539230 582648
rect 480200 573864 496200 581588
rect 516200 581478 539230 582014
rect 523230 573830 539230 581478
rect 30318 561264 46318 569418
rect 57044 568200 58054 568400
rect 57044 567720 57198 568200
rect 57918 567720 58054 568200
rect 57044 567300 58054 567720
rect 60764 568200 61774 568400
rect 60764 567720 60918 568200
rect 61638 567720 61774 568200
rect 57064 561264 58032 567300
rect 60764 561428 61774 567720
rect 60730 561412 63776 561428
rect 73428 561412 89428 569276
rect 30318 560338 58072 561264
rect 30318 553218 46318 560338
rect 60730 560296 89428 561412
rect 73400 560188 89428 560296
rect 73428 553076 89428 560188
rect 120318 561264 136318 569418
rect 147044 568200 148054 568400
rect 147044 567720 147198 568200
rect 147918 567720 148054 568200
rect 147044 567300 148054 567720
rect 150764 568200 151774 568400
rect 150764 567720 150918 568200
rect 151638 567720 151774 568200
rect 147064 561264 148032 567300
rect 150764 561428 151774 567720
rect 150730 561412 153776 561428
rect 163428 561412 179428 569276
rect 120318 560338 148072 561264
rect 120318 553218 136318 560338
rect 150730 560296 179428 561412
rect 163400 560188 179428 560296
rect 163428 553076 179428 560188
rect 210318 561264 226318 569418
rect 237044 568200 238054 568400
rect 237044 567720 237198 568200
rect 237918 567720 238054 568200
rect 237044 567300 238054 567720
rect 240764 568200 241774 568400
rect 240764 567720 240918 568200
rect 241638 567720 241774 568200
rect 237064 561264 238032 567300
rect 240764 561428 241774 567720
rect 240730 561412 243776 561428
rect 253428 561412 269428 569276
rect 210318 560338 238072 561264
rect 210318 553218 226318 560338
rect 240730 560296 269428 561412
rect 253400 560188 269428 560296
rect 253428 553076 269428 560188
rect 300318 561264 316318 569418
rect 327044 568200 328054 568400
rect 327044 567720 327198 568200
rect 327918 567720 328054 568200
rect 327044 567300 328054 567720
rect 330764 568200 331774 568400
rect 330764 567720 330918 568200
rect 331638 567720 331774 568200
rect 327064 561264 328032 567300
rect 330764 561428 331774 567720
rect 330730 561412 333776 561428
rect 343428 561412 359428 569276
rect 300318 560338 328072 561264
rect 300318 553218 316318 560338
rect 330730 560296 359428 561412
rect 343400 560188 359428 560296
rect 343428 553076 359428 560188
rect 390120 563188 406120 571342
rect 416846 570124 417856 570324
rect 416846 569644 417000 570124
rect 417720 569644 417856 570124
rect 416846 569224 417856 569644
rect 420566 570124 421576 570324
rect 420566 569644 420720 570124
rect 421440 569644 421576 570124
rect 416866 563188 417834 569224
rect 420566 563352 421576 569644
rect 420532 563336 423578 563352
rect 433230 563336 449230 571200
rect 390120 562262 417874 563188
rect 390120 555142 406120 562262
rect 420532 562220 449230 563336
rect 433202 562112 449230 562220
rect 433230 555000 449230 562112
rect 480120 563188 496120 571342
rect 506846 570124 507856 570324
rect 506846 569644 507000 570124
rect 507720 569644 507856 570124
rect 506846 569224 507856 569644
rect 510566 570124 511576 570324
rect 510566 569644 510720 570124
rect 511440 569644 511576 570124
rect 506866 563188 507834 569224
rect 510566 563352 511576 569644
rect 510532 563336 513578 563352
rect 523230 563336 539230 571200
rect 480120 562262 507874 563188
rect 480120 555142 496120 562262
rect 510532 562220 539230 563336
rect 523202 562112 539230 562220
rect 523230 555000 539230 562112
rect 51294 517964 67294 534164
rect 141294 517964 157294 534164
rect 231294 517964 247294 534164
rect 321294 517964 337294 534164
rect 411294 517964 427294 534164
rect 501294 517964 517294 534164
rect 30332 512300 46332 517920
rect 63816 516794 66376 517964
rect 63816 515116 64332 516794
rect 65752 515116 66376 516794
rect 63816 514208 66376 515116
rect 30332 511040 58098 512300
rect 73518 512240 89518 517940
rect 72558 512224 89518 512240
rect 60790 511108 89518 512224
rect 60790 511092 63836 511108
rect 72558 511100 89518 511108
rect 30332 509140 46332 511040
rect 30198 508140 46338 509140
rect 30332 501720 46332 508140
rect 57124 505220 58092 511040
rect 57104 504800 58114 505220
rect 57104 504320 57258 504800
rect 57978 504320 58114 504800
rect 57104 504120 58114 504320
rect 60824 504800 61834 511092
rect 60824 504320 60978 504800
rect 61698 504320 61834 504800
rect 60824 504120 61834 504320
rect 73518 501740 89518 511100
rect 120332 512300 136332 517920
rect 153816 516794 156376 517964
rect 153816 515116 154332 516794
rect 155752 515116 156376 516794
rect 153816 514208 156376 515116
rect 120332 511040 148098 512300
rect 163518 512240 179518 517940
rect 162558 512224 179518 512240
rect 150790 511108 179518 512224
rect 150790 511092 153836 511108
rect 162558 511100 179518 511108
rect 120332 509140 136332 511040
rect 120198 508140 136338 509140
rect 120332 501720 136332 508140
rect 147124 505220 148092 511040
rect 147104 504800 148114 505220
rect 147104 504320 147258 504800
rect 147978 504320 148114 504800
rect 147104 504120 148114 504320
rect 150824 504800 151834 511092
rect 150824 504320 150978 504800
rect 151698 504320 151834 504800
rect 150824 504120 151834 504320
rect 163518 501740 179518 511100
rect 210332 512300 226332 517920
rect 243816 516794 246376 517964
rect 243816 515116 244332 516794
rect 245752 515116 246376 516794
rect 243816 514208 246376 515116
rect 210332 511040 238098 512300
rect 253518 512240 269518 517940
rect 252558 512224 269518 512240
rect 240790 511108 269518 512224
rect 240790 511092 243836 511108
rect 252558 511100 269518 511108
rect 210332 509140 226332 511040
rect 210198 508140 226338 509140
rect 210332 501720 226332 508140
rect 237124 505220 238092 511040
rect 237104 504800 238114 505220
rect 237104 504320 237258 504800
rect 237978 504320 238114 504800
rect 237104 504120 238114 504320
rect 240824 504800 241834 511092
rect 240824 504320 240978 504800
rect 241698 504320 241834 504800
rect 240824 504120 241834 504320
rect 253518 501740 269518 511100
rect 300332 512300 316332 517920
rect 333816 516794 336376 517964
rect 333816 515116 334332 516794
rect 335752 515116 336376 516794
rect 333816 514208 336376 515116
rect 300332 511040 328098 512300
rect 343518 512240 359518 517940
rect 342558 512224 359518 512240
rect 330790 511108 359518 512224
rect 330790 511092 333836 511108
rect 342558 511100 359518 511108
rect 300332 509140 316332 511040
rect 300198 508140 316338 509140
rect 300332 501720 316332 508140
rect 327124 505220 328092 511040
rect 327104 504800 328114 505220
rect 327104 504320 327258 504800
rect 327978 504320 328114 504800
rect 327104 504120 328114 504320
rect 330824 504800 331834 511092
rect 330824 504320 330978 504800
rect 331698 504320 331834 504800
rect 330824 504120 331834 504320
rect 343518 501740 359518 511100
rect 390332 512300 406332 517920
rect 423816 516794 426376 517964
rect 423816 515116 424332 516794
rect 425752 515116 426376 516794
rect 423816 514208 426376 515116
rect 390332 511040 418098 512300
rect 433518 512240 449518 517940
rect 432558 512224 449518 512240
rect 420790 511108 449518 512224
rect 420790 511092 423836 511108
rect 432558 511100 449518 511108
rect 390332 509140 406332 511040
rect 390198 508140 406338 509140
rect 390332 501720 406332 508140
rect 417124 505220 418092 511040
rect 417104 504800 418114 505220
rect 417104 504320 417258 504800
rect 417978 504320 418114 504800
rect 417104 504120 418114 504320
rect 420824 504800 421834 511092
rect 420824 504320 420978 504800
rect 421698 504320 421834 504800
rect 420824 504120 421834 504320
rect 433518 501740 449518 511100
rect 480332 512300 496332 517920
rect 513816 516794 516376 517964
rect 513816 515116 514332 516794
rect 515752 515116 516376 516794
rect 513816 514208 516376 515116
rect 480332 511040 508098 512300
rect 523518 512240 539518 517940
rect 522558 512224 539518 512240
rect 510790 511108 539518 512224
rect 510790 511092 513836 511108
rect 522558 511100 539518 511108
rect 480332 509140 496332 511040
rect 480198 508140 496338 509140
rect 480332 501720 496332 508140
rect 507124 505220 508092 511040
rect 507104 504800 508114 505220
rect 507104 504320 507258 504800
rect 507978 504320 508114 504800
rect 507104 504120 508114 504320
rect 510824 504800 511834 511092
rect 510824 504320 510978 504800
rect 511698 504320 511834 504800
rect 510824 504120 511834 504320
rect 523518 501740 539518 511100
rect 30398 492054 46398 499240
rect 73428 492194 89428 499206
rect 30398 492050 53488 492054
rect 30398 491360 53546 492050
rect 30398 491040 53194 491360
rect 53514 491040 53546 491360
rect 30398 490764 53546 491040
rect 66398 491824 89428 492194
rect 66398 491190 66566 491824
rect 67218 491190 89428 491824
rect 30398 483040 46398 490764
rect 66398 490654 89428 491190
rect 73428 483006 89428 490654
rect 120398 492054 136398 499240
rect 163428 492194 179428 499206
rect 120398 490764 136428 492054
rect 120398 485900 136398 490764
rect 163413 490654 179428 492194
rect 160159 487410 161077 487434
rect 163428 487410 179428 490654
rect 160159 486540 160183 487410
rect 161053 486540 179428 487410
rect 160159 486516 161077 486540
rect 139639 485900 140777 485924
rect 120398 484810 139663 485900
rect 140753 484810 140777 485900
rect 120398 483040 136398 484810
rect 139639 484786 140777 484810
rect 163428 483006 179428 486540
rect 210398 492054 226398 499240
rect 253428 492194 269428 499206
rect 249801 492164 251350 492187
rect 252749 492164 269428 492194
rect 249801 492163 269428 492164
rect 210398 491779 226416 492054
rect 210398 491774 226774 491779
rect 227645 491774 228641 491798
rect 210398 490826 227669 491774
rect 228617 490826 228641 491774
rect 210398 490825 226774 490826
rect 210398 490764 226402 490825
rect 227645 490802 228641 490826
rect 210398 483040 226398 490764
rect 249801 490662 249825 492163
rect 251326 490663 269428 492163
rect 251326 490662 251350 490663
rect 249801 490638 251350 490662
rect 252749 490654 269428 490663
rect 253428 483006 269428 490654
rect 300398 492054 316398 499240
rect 343428 492194 359428 499206
rect 300398 491749 318624 492054
rect 319603 491749 319977 491773
rect 300398 491423 319627 491749
rect 319953 491423 319977 491749
rect 300398 490764 318624 491423
rect 319603 491399 319977 491423
rect 341132 491700 359428 492194
rect 341132 491278 341405 491700
rect 341827 491278 359428 491700
rect 300398 483040 316398 490764
rect 341132 490654 359428 491278
rect 343428 483006 359428 490654
rect 390398 492054 406398 499240
rect 433428 492194 449428 499206
rect 390398 492050 413488 492054
rect 390398 491360 413546 492050
rect 390398 491040 413194 491360
rect 413514 491040 413546 491360
rect 390398 490764 413546 491040
rect 426398 491824 449428 492194
rect 426398 491190 426566 491824
rect 427218 491190 449428 491824
rect 390398 483040 406398 490764
rect 426398 490654 449428 491190
rect 433428 483006 449428 490654
rect 480398 492054 496398 499240
rect 523428 492194 539428 499206
rect 480398 492050 503488 492054
rect 480398 491360 503546 492050
rect 480398 491040 503194 491360
rect 503514 491040 503546 491360
rect 480398 490764 503546 491040
rect 516398 491824 539428 492194
rect 516398 491190 516566 491824
rect 517218 491190 539428 491824
rect 480398 483040 496398 490764
rect 516398 490654 539428 491190
rect 523428 483006 539428 490654
rect 30318 472364 46318 480518
rect 57044 479300 58054 479500
rect 57044 478820 57198 479300
rect 57918 478820 58054 479300
rect 57044 478400 58054 478820
rect 60764 479300 61774 479500
rect 60764 478820 60918 479300
rect 61638 478820 61774 479300
rect 57064 472364 58032 478400
rect 60764 472528 61774 478820
rect 60730 472512 63776 472528
rect 73428 472512 89428 480376
rect 30318 471438 58072 472364
rect 30318 464318 46318 471438
rect 60730 471396 89428 472512
rect 73400 471288 89428 471396
rect 51806 468222 54366 469006
rect 51806 466544 52334 468222
rect 53754 466544 54366 468222
rect 51806 464276 54366 466544
rect 50782 448076 66782 464276
rect 73428 464176 89428 471288
rect 120318 472364 136318 480518
rect 147044 479300 148054 479500
rect 147044 478820 147198 479300
rect 147918 478820 148054 479300
rect 147044 478400 148054 478820
rect 150764 479300 151774 479500
rect 150764 478820 150918 479300
rect 151638 478820 151774 479300
rect 147064 472364 148032 478400
rect 150764 472528 151774 478820
rect 150730 472512 153776 472528
rect 163428 472512 179428 480376
rect 120318 471438 148072 472364
rect 120318 464318 136318 471438
rect 150730 471396 179428 472512
rect 163400 471288 179428 471396
rect 141806 468222 144366 469006
rect 141806 466544 142334 468222
rect 143754 466544 144366 468222
rect 141806 464276 144366 466544
rect 140782 448076 156782 464276
rect 163428 464176 179428 471288
rect 210318 472364 226318 480518
rect 237044 479300 238054 479500
rect 237044 478820 237198 479300
rect 237918 478820 238054 479300
rect 237044 478400 238054 478820
rect 240764 479300 241774 479500
rect 240764 478820 240918 479300
rect 241638 478820 241774 479300
rect 237064 472364 238032 478400
rect 240764 472528 241774 478820
rect 240730 472512 243776 472528
rect 253428 472512 269428 480376
rect 210318 471438 238072 472364
rect 210318 464318 226318 471438
rect 240730 471396 269428 472512
rect 253400 471288 269428 471396
rect 231806 468222 234366 469006
rect 231806 466544 232334 468222
rect 233754 466544 234366 468222
rect 231806 464276 234366 466544
rect 230782 448076 246782 464276
rect 253428 464176 269428 471288
rect 300318 472364 316318 480518
rect 327044 479300 328054 479500
rect 327044 478820 327198 479300
rect 327918 478820 328054 479300
rect 327044 478400 328054 478820
rect 330764 479300 331774 479500
rect 330764 478820 330918 479300
rect 331638 478820 331774 479300
rect 327064 472364 328032 478400
rect 330764 472528 331774 478820
rect 330730 472512 333776 472528
rect 343428 472512 359428 480376
rect 300318 471438 328072 472364
rect 300318 464318 316318 471438
rect 330730 471396 359428 472512
rect 343400 471288 359428 471396
rect 321806 468222 324366 469006
rect 321806 466544 322334 468222
rect 323754 466544 324366 468222
rect 321806 464276 324366 466544
rect 320782 448076 336782 464276
rect 343428 464176 359428 471288
rect 390318 472364 406318 480518
rect 417044 479300 418054 479500
rect 417044 478820 417198 479300
rect 417918 478820 418054 479300
rect 417044 478400 418054 478820
rect 420764 479300 421774 479500
rect 420764 478820 420918 479300
rect 421638 478820 421774 479300
rect 417064 472364 418032 478400
rect 420764 472528 421774 478820
rect 420730 472512 423776 472528
rect 433428 472512 449428 480376
rect 390318 471438 418072 472364
rect 390318 464318 406318 471438
rect 420730 471396 449428 472512
rect 433400 471288 449428 471396
rect 411806 468222 414366 469006
rect 411806 466544 412334 468222
rect 413754 466544 414366 468222
rect 411806 464276 414366 466544
rect 410782 448076 426782 464276
rect 433428 464176 449428 471288
rect 480318 472364 496318 480518
rect 507044 479300 508054 479500
rect 507044 478820 507198 479300
rect 507918 478820 508054 479300
rect 507044 478400 508054 478820
rect 510764 479300 511774 479500
rect 510764 478820 510918 479300
rect 511638 478820 511774 479300
rect 507064 472364 508032 478400
rect 510764 472528 511774 478820
rect 510730 472512 513776 472528
rect 523428 472512 539428 480376
rect 480318 471438 508072 472364
rect 480318 464318 496318 471438
rect 510730 471396 539428 472512
rect 523400 471288 539428 471396
rect 501806 468222 504366 469006
rect 501806 466544 502334 468222
rect 503754 466544 504366 468222
rect 501806 464276 504366 466544
rect 500782 448076 516782 464276
rect 523428 464176 539428 471288
rect 51294 397964 67294 414164
rect 141294 397964 157294 414164
rect 231294 397964 247294 414164
rect 321294 397964 337294 414164
rect 411294 397964 427294 414164
rect 501294 397964 517294 414164
rect 30332 392300 46332 397920
rect 63816 396794 66376 397964
rect 63816 395116 64332 396794
rect 65752 395116 66376 396794
rect 63816 394208 66376 395116
rect 30332 391040 58098 392300
rect 73518 392240 89518 397940
rect 72558 392224 89518 392240
rect 60790 391108 89518 392224
rect 60790 391092 63836 391108
rect 72558 391100 89518 391108
rect 30332 389140 46332 391040
rect 30198 388140 46338 389140
rect 30332 381720 46332 388140
rect 57124 385220 58092 391040
rect 57104 384800 58114 385220
rect 57104 384320 57258 384800
rect 57978 384320 58114 384800
rect 57104 384120 58114 384320
rect 60824 384800 61834 391092
rect 60824 384320 60978 384800
rect 61698 384320 61834 384800
rect 60824 384120 61834 384320
rect 73518 381740 89518 391100
rect 120332 392300 136332 397920
rect 153816 396794 156376 397964
rect 153816 395116 154332 396794
rect 155752 395116 156376 396794
rect 153816 394208 156376 395116
rect 120332 391040 148098 392300
rect 163518 392240 179518 397940
rect 162558 392224 179518 392240
rect 150790 391108 179518 392224
rect 150790 391092 153836 391108
rect 162558 391100 179518 391108
rect 120332 389140 136332 391040
rect 120198 388140 136338 389140
rect 120332 381720 136332 388140
rect 147124 385220 148092 391040
rect 147104 384800 148114 385220
rect 147104 384320 147258 384800
rect 147978 384320 148114 384800
rect 147104 384120 148114 384320
rect 150824 384800 151834 391092
rect 150824 384320 150978 384800
rect 151698 384320 151834 384800
rect 150824 384120 151834 384320
rect 163518 381740 179518 391100
rect 210332 392300 226332 397920
rect 243816 396794 246376 397964
rect 243816 395116 244332 396794
rect 245752 395116 246376 396794
rect 243816 394208 246376 395116
rect 210332 391040 238098 392300
rect 253518 392240 269518 397940
rect 252558 392224 269518 392240
rect 240790 391108 269518 392224
rect 240790 391092 243836 391108
rect 252558 391100 269518 391108
rect 210332 389140 226332 391040
rect 210198 388140 226338 389140
rect 210332 381720 226332 388140
rect 237124 385220 238092 391040
rect 237104 384800 238114 385220
rect 237104 384320 237258 384800
rect 237978 384320 238114 384800
rect 237104 384120 238114 384320
rect 240824 384800 241834 391092
rect 240824 384320 240978 384800
rect 241698 384320 241834 384800
rect 240824 384120 241834 384320
rect 253518 381740 269518 391100
rect 300332 392300 316332 397920
rect 333816 396794 336376 397964
rect 333816 395116 334332 396794
rect 335752 395116 336376 396794
rect 333816 394208 336376 395116
rect 300332 391040 328098 392300
rect 343518 392240 359518 397940
rect 342558 392224 359518 392240
rect 330790 391108 359518 392224
rect 330790 391092 333836 391108
rect 342558 391100 359518 391108
rect 300332 389140 316332 391040
rect 300198 388140 316338 389140
rect 300332 381720 316332 388140
rect 327124 385220 328092 391040
rect 327104 384800 328114 385220
rect 327104 384320 327258 384800
rect 327978 384320 328114 384800
rect 327104 384120 328114 384320
rect 330824 384800 331834 391092
rect 330824 384320 330978 384800
rect 331698 384320 331834 384800
rect 330824 384120 331834 384320
rect 343518 381740 359518 391100
rect 390332 392300 406332 397920
rect 423816 396794 426376 397964
rect 423816 395116 424332 396794
rect 425752 395116 426376 396794
rect 423816 394208 426376 395116
rect 390332 391040 418098 392300
rect 433518 392240 449518 397940
rect 432558 392224 449518 392240
rect 420790 391108 449518 392224
rect 420790 391092 423836 391108
rect 432558 391100 449518 391108
rect 390332 389140 406332 391040
rect 390198 388140 406338 389140
rect 390332 381720 406332 388140
rect 417124 385220 418092 391040
rect 417104 384800 418114 385220
rect 417104 384320 417258 384800
rect 417978 384320 418114 384800
rect 417104 384120 418114 384320
rect 420824 384800 421834 391092
rect 420824 384320 420978 384800
rect 421698 384320 421834 384800
rect 420824 384120 421834 384320
rect 433518 381740 449518 391100
rect 480332 392300 496332 397920
rect 513816 396794 516376 397964
rect 513816 395116 514332 396794
rect 515752 395116 516376 396794
rect 513816 394208 516376 395116
rect 480332 391040 508098 392300
rect 523518 392240 539518 397940
rect 522558 392224 539518 392240
rect 510790 391108 539518 392224
rect 510790 391092 513836 391108
rect 522558 391100 539518 391108
rect 480332 389140 496332 391040
rect 480198 388140 496338 389140
rect 480332 381720 496332 388140
rect 507124 385220 508092 391040
rect 507104 384800 508114 385220
rect 507104 384320 507258 384800
rect 507978 384320 508114 384800
rect 507104 384120 508114 384320
rect 510824 384800 511834 391092
rect 510824 384320 510978 384800
rect 511698 384320 511834 384800
rect 510824 384120 511834 384320
rect 523518 381740 539518 391100
rect 30398 372054 46398 379240
rect 73428 372194 89428 379206
rect 30398 370764 46428 372054
rect 30398 365900 46398 370764
rect 73413 370654 89428 372194
rect 70159 367410 71077 367434
rect 73428 367410 89428 370654
rect 70159 366540 70183 367410
rect 71053 366540 89428 367410
rect 70159 366516 71077 366540
rect 49639 365900 50777 365924
rect 30398 364810 49663 365900
rect 50753 364810 50777 365900
rect 30398 363040 46398 364810
rect 49639 364786 50777 364810
rect 73428 363006 89428 366540
rect 120398 372054 136398 379240
rect 163428 372194 179428 379206
rect 120398 370764 136428 372054
rect 120398 365900 136398 370764
rect 163413 370654 179428 372194
rect 160159 367410 161077 367434
rect 163428 367410 179428 370654
rect 160159 366540 160183 367410
rect 161053 366540 179428 367410
rect 160159 366516 161077 366540
rect 139639 365900 140777 365924
rect 120398 364810 139663 365900
rect 140753 364810 140777 365900
rect 120398 363040 136398 364810
rect 139639 364786 140777 364810
rect 163428 363006 179428 366540
rect 210398 372054 226398 379240
rect 253428 372194 269428 379206
rect 249801 372164 251350 372187
rect 252749 372164 269428 372194
rect 249801 372163 269428 372164
rect 210398 371779 226416 372054
rect 210398 371774 226774 371779
rect 227645 371774 228641 371798
rect 210398 370826 227669 371774
rect 228617 370826 228641 371774
rect 210398 370825 226774 370826
rect 210398 370764 226402 370825
rect 227645 370802 228641 370826
rect 210398 363040 226398 370764
rect 249801 370662 249825 372163
rect 251326 370663 269428 372163
rect 251326 370662 251350 370663
rect 249801 370638 251350 370662
rect 252749 370654 269428 370663
rect 253428 363006 269428 370654
rect 300398 372054 316398 379240
rect 343428 372194 359428 379206
rect 300398 371749 318624 372054
rect 319603 371749 319977 371773
rect 300398 371423 319627 371749
rect 319953 371423 319977 371749
rect 300398 370764 318624 371423
rect 319603 371399 319977 371423
rect 341132 371700 359428 372194
rect 341132 371278 341405 371700
rect 341827 371278 359428 371700
rect 300398 363040 316398 370764
rect 341132 370654 359428 371278
rect 343428 363006 359428 370654
rect 390398 372054 406398 379240
rect 433428 372194 449428 379206
rect 390398 372050 413488 372054
rect 390398 371360 413546 372050
rect 390398 371040 413194 371360
rect 413514 371040 413546 371360
rect 390398 370764 413546 371040
rect 426398 371824 449428 372194
rect 426398 371190 426566 371824
rect 427218 371190 449428 371824
rect 390398 363040 406398 370764
rect 426398 370654 449428 371190
rect 433428 363006 449428 370654
rect 480398 372054 496398 379240
rect 523428 372194 539428 379206
rect 480398 372050 503488 372054
rect 480398 371360 503546 372050
rect 480398 371040 503194 371360
rect 503514 371040 503546 371360
rect 480398 370764 503546 371040
rect 516398 371824 539428 372194
rect 516398 371190 516566 371824
rect 517218 371190 539428 371824
rect 480398 363040 496398 370764
rect 516398 370654 539428 371190
rect 523428 363006 539428 370654
rect 30318 352364 46318 360518
rect 57044 359300 58054 359500
rect 57044 358820 57198 359300
rect 57918 358820 58054 359300
rect 57044 358400 58054 358820
rect 60764 359300 61774 359500
rect 60764 358820 60918 359300
rect 61638 358820 61774 359300
rect 57064 352364 58032 358400
rect 60764 352528 61774 358820
rect 60730 352512 63776 352528
rect 73428 352512 89428 360376
rect 30318 351438 58072 352364
rect 30318 344318 46318 351438
rect 60730 351396 89428 352512
rect 73400 351288 89428 351396
rect 51806 348222 54366 349006
rect 51806 346544 52334 348222
rect 53754 346544 54366 348222
rect 51806 344276 54366 346544
rect 50782 328076 66782 344276
rect 73428 344176 89428 351288
rect 120318 352364 136318 360518
rect 147044 359300 148054 359500
rect 147044 358820 147198 359300
rect 147918 358820 148054 359300
rect 147044 358400 148054 358820
rect 150764 359300 151774 359500
rect 150764 358820 150918 359300
rect 151638 358820 151774 359300
rect 147064 352364 148032 358400
rect 150764 352528 151774 358820
rect 150730 352512 153776 352528
rect 163428 352512 179428 360376
rect 120318 351438 148072 352364
rect 120318 344318 136318 351438
rect 150730 351396 179428 352512
rect 163400 351288 179428 351396
rect 141806 348222 144366 349006
rect 141806 346544 142334 348222
rect 143754 346544 144366 348222
rect 141806 344276 144366 346544
rect 140782 328076 156782 344276
rect 163428 344176 179428 351288
rect 210318 352364 226318 360518
rect 237044 359300 238054 359500
rect 237044 358820 237198 359300
rect 237918 358820 238054 359300
rect 237044 358400 238054 358820
rect 240764 359300 241774 359500
rect 240764 358820 240918 359300
rect 241638 358820 241774 359300
rect 237064 352364 238032 358400
rect 240764 352528 241774 358820
rect 240730 352512 243776 352528
rect 253428 352512 269428 360376
rect 210318 351438 238072 352364
rect 210318 344318 226318 351438
rect 240730 351396 269428 352512
rect 253400 351288 269428 351396
rect 231806 348222 234366 349006
rect 231806 346544 232334 348222
rect 233754 346544 234366 348222
rect 231806 344276 234366 346544
rect 230782 328076 246782 344276
rect 253428 344176 269428 351288
rect 300318 352364 316318 360518
rect 327044 359300 328054 359500
rect 327044 358820 327198 359300
rect 327918 358820 328054 359300
rect 327044 358400 328054 358820
rect 330764 359300 331774 359500
rect 330764 358820 330918 359300
rect 331638 358820 331774 359300
rect 327064 352364 328032 358400
rect 330764 352528 331774 358820
rect 330730 352512 333776 352528
rect 343428 352512 359428 360376
rect 300318 351438 328072 352364
rect 300318 344318 316318 351438
rect 330730 351396 359428 352512
rect 343400 351288 359428 351396
rect 321806 348222 324366 349006
rect 321806 346544 322334 348222
rect 323754 346544 324366 348222
rect 321806 344276 324366 346544
rect 320782 328076 336782 344276
rect 343428 344176 359428 351288
rect 390318 352364 406318 360518
rect 417044 359300 418054 359500
rect 417044 358820 417198 359300
rect 417918 358820 418054 359300
rect 417044 358400 418054 358820
rect 420764 359300 421774 359500
rect 420764 358820 420918 359300
rect 421638 358820 421774 359300
rect 417064 352364 418032 358400
rect 420764 352528 421774 358820
rect 420730 352512 423776 352528
rect 433428 352512 449428 360376
rect 390318 351438 418072 352364
rect 390318 344318 406318 351438
rect 420730 351396 449428 352512
rect 433400 351288 449428 351396
rect 411806 348222 414366 349006
rect 411806 346544 412334 348222
rect 413754 346544 414366 348222
rect 411806 344276 414366 346544
rect 410782 328076 426782 344276
rect 433428 344176 449428 351288
rect 480318 352364 496318 360518
rect 507044 359300 508054 359500
rect 507044 358820 507198 359300
rect 507918 358820 508054 359300
rect 507044 358400 508054 358820
rect 510764 359300 511774 359500
rect 510764 358820 510918 359300
rect 511638 358820 511774 359300
rect 507064 352364 508032 358400
rect 510764 352528 511774 358820
rect 510730 352512 513776 352528
rect 523428 352512 539428 360376
rect 480318 351438 508072 352364
rect 480318 344318 496318 351438
rect 510730 351396 539428 352512
rect 523400 351288 539428 351396
rect 501806 348222 504366 349006
rect 501806 346544 502334 348222
rect 503754 346544 504366 348222
rect 501806 344276 504366 346544
rect 500782 328076 516782 344276
rect 523428 344176 539428 351288
rect 51294 277964 67294 294164
rect 30332 272300 46332 277920
rect 63816 276794 66376 277964
rect 63816 275116 64332 276794
rect 65752 275116 66376 276794
rect 63816 274208 66376 275116
rect 30332 271040 58098 272300
rect 73518 272240 89518 277940
rect 140418 277760 156418 293960
rect 72558 272224 89518 272240
rect 60790 271108 89518 272224
rect 60790 271092 63836 271108
rect 72558 271100 89518 271108
rect 30332 269140 46332 271040
rect 30198 268140 46338 269140
rect 30332 261720 46332 268140
rect 57124 265220 58092 271040
rect 57104 264800 58114 265220
rect 57104 264320 57258 264800
rect 57978 264320 58114 264800
rect 57104 264120 58114 264320
rect 60824 264800 61834 271092
rect 60824 264320 60978 264800
rect 61698 264320 61834 264800
rect 60824 264120 61834 264320
rect 73518 261740 89518 271100
rect 119456 272096 135456 277716
rect 152940 276590 155500 277760
rect 152940 274912 153456 276590
rect 154876 274912 155500 276590
rect 152940 274004 155500 274912
rect 119456 270836 147222 272096
rect 162642 272036 178642 277736
rect 231672 277572 247672 293772
rect 321294 277964 337294 294164
rect 411294 277964 427294 294164
rect 501294 277964 517294 294164
rect 161682 272020 178642 272036
rect 149914 270904 178642 272020
rect 149914 270888 152960 270904
rect 161682 270896 178642 270904
rect 119456 268936 135456 270836
rect 119322 267936 135462 268936
rect 119456 261516 135456 267936
rect 146248 265016 147216 270836
rect 146228 264596 147238 265016
rect 146228 264116 146382 264596
rect 147102 264116 147238 264596
rect 146228 263916 147238 264116
rect 149948 264596 150958 270888
rect 149948 264116 150102 264596
rect 150822 264116 150958 264596
rect 149948 263916 150958 264116
rect 162642 261536 178642 270896
rect 210710 271908 226710 277528
rect 244194 276402 246754 277572
rect 244194 274724 244710 276402
rect 246130 274724 246754 276402
rect 244194 273816 246754 274724
rect 210710 270648 238476 271908
rect 253896 271848 269896 277548
rect 252936 271832 269896 271848
rect 241168 270716 269896 271832
rect 241168 270700 244214 270716
rect 252936 270708 269896 270716
rect 210710 268748 226710 270648
rect 210576 267748 226716 268748
rect 210710 261328 226710 267748
rect 237502 264828 238470 270648
rect 237482 264408 238492 264828
rect 237482 263928 237636 264408
rect 238356 263928 238492 264408
rect 237482 263728 238492 263928
rect 241202 264408 242212 270700
rect 241202 263928 241356 264408
rect 242076 263928 242212 264408
rect 241202 263728 242212 263928
rect 253896 261348 269896 270708
rect 300332 272300 316332 277920
rect 333816 276794 336376 277964
rect 333816 275116 334332 276794
rect 335752 275116 336376 276794
rect 333816 274208 336376 275116
rect 300332 271040 328098 272300
rect 343518 272240 359518 277940
rect 342558 272224 359518 272240
rect 330790 271108 359518 272224
rect 330790 271092 333836 271108
rect 342558 271100 359518 271108
rect 300332 269140 316332 271040
rect 300198 268140 316338 269140
rect 300332 261720 316332 268140
rect 327124 265220 328092 271040
rect 327104 264800 328114 265220
rect 327104 264320 327258 264800
rect 327978 264320 328114 264800
rect 327104 264120 328114 264320
rect 330824 264800 331834 271092
rect 330824 264320 330978 264800
rect 331698 264320 331834 264800
rect 330824 264120 331834 264320
rect 343518 261740 359518 271100
rect 390332 272300 406332 277920
rect 423816 276794 426376 277964
rect 423816 275116 424332 276794
rect 425752 275116 426376 276794
rect 423816 274208 426376 275116
rect 390332 271040 418098 272300
rect 433518 272240 449518 277940
rect 432558 272224 449518 272240
rect 420790 271108 449518 272224
rect 420790 271092 423836 271108
rect 432558 271100 449518 271108
rect 390332 269140 406332 271040
rect 390198 268140 406338 269140
rect 390332 261720 406332 268140
rect 417124 265220 418092 271040
rect 417104 264800 418114 265220
rect 417104 264320 417258 264800
rect 417978 264320 418114 264800
rect 417104 264120 418114 264320
rect 420824 264800 421834 271092
rect 420824 264320 420978 264800
rect 421698 264320 421834 264800
rect 420824 264120 421834 264320
rect 433518 261740 449518 271100
rect 480332 272300 496332 277920
rect 513816 276794 516376 277964
rect 513816 275116 514332 276794
rect 515752 275116 516376 276794
rect 513816 274208 516376 275116
rect 480332 271040 508098 272300
rect 523518 272240 539518 277940
rect 522558 272224 539518 272240
rect 510790 271108 539518 272224
rect 510790 271092 513836 271108
rect 522558 271100 539518 271108
rect 480332 269140 496332 271040
rect 480198 268140 496338 269140
rect 480332 261720 496332 268140
rect 507124 265220 508092 271040
rect 507104 264800 508114 265220
rect 507104 264320 507258 264800
rect 507978 264320 508114 264800
rect 507104 264120 508114 264320
rect 510824 264800 511834 271092
rect 510824 264320 510978 264800
rect 511698 264320 511834 264800
rect 510824 264120 511834 264320
rect 523518 261740 539518 271100
rect 30398 252054 46398 259240
rect 73428 252194 89428 259206
rect 30398 252050 53488 252054
rect 30398 251360 53546 252050
rect 30398 251040 53194 251360
rect 53514 251040 53546 251360
rect 30398 250764 53546 251040
rect 66398 251824 89428 252194
rect 66398 251190 66566 251824
rect 67218 251190 89428 251824
rect 30398 243040 46398 250764
rect 66398 250654 89428 251190
rect 73428 243006 89428 250654
rect 119522 251850 135522 259036
rect 162552 251990 178552 259002
rect 119522 251846 142612 251850
rect 119522 251156 142670 251846
rect 119522 250836 142318 251156
rect 142638 250836 142670 251156
rect 119522 250560 142670 250836
rect 155522 251620 178552 251990
rect 155522 250986 155690 251620
rect 156342 250986 178552 251620
rect 119522 242836 135522 250560
rect 155522 250450 178552 250986
rect 162552 242802 178552 250450
rect 210776 251662 226776 258848
rect 253806 251802 269806 258814
rect 210776 251357 229002 251662
rect 229981 251357 230355 251381
rect 210776 251031 230005 251357
rect 230331 251031 230355 251357
rect 210776 250372 229002 251031
rect 229981 251007 230355 251031
rect 251510 251308 269806 251802
rect 251510 250886 251783 251308
rect 252205 250886 269806 251308
rect 210776 242648 226776 250372
rect 251510 250262 269806 250886
rect 253806 242614 269806 250262
rect 300398 252054 316398 259240
rect 343428 252194 359428 259206
rect 339801 252164 341350 252187
rect 342749 252164 359428 252194
rect 339801 252163 359428 252164
rect 300398 251779 316416 252054
rect 300398 251774 316774 251779
rect 317645 251774 318641 251798
rect 300398 250826 317669 251774
rect 318617 250826 318641 251774
rect 300398 250825 316774 250826
rect 300398 250764 316402 250825
rect 317645 250802 318641 250826
rect 300398 243040 316398 250764
rect 339801 250662 339825 252163
rect 341326 250663 359428 252163
rect 341326 250662 341350 250663
rect 339801 250638 341350 250662
rect 342749 250654 359428 250663
rect 343428 243006 359428 250654
rect 390398 252054 406398 259240
rect 433428 252194 449428 259206
rect 390398 250764 406428 252054
rect 390398 245900 406398 250764
rect 433413 250654 449428 252194
rect 430159 247410 431077 247434
rect 433428 247410 449428 250654
rect 430159 246540 430183 247410
rect 431053 246540 449428 247410
rect 430159 246516 431077 246540
rect 409639 245900 410777 245924
rect 390398 244810 409663 245900
rect 410753 244810 410777 245900
rect 390398 243040 406398 244810
rect 409639 244786 410777 244810
rect 433428 243006 449428 246540
rect 480398 252054 496398 259240
rect 523428 252194 539428 259206
rect 480398 250764 496428 252054
rect 480398 245900 496398 250764
rect 523413 250654 539428 252194
rect 520159 247410 521077 247434
rect 523428 247410 539428 250654
rect 520159 246540 520183 247410
rect 521053 246540 539428 247410
rect 520159 246516 521077 246540
rect 499639 245900 500777 245924
rect 480398 244810 499663 245900
rect 500753 244810 500777 245900
rect 480398 243040 496398 244810
rect 499639 244786 500777 244810
rect 523428 243006 539428 246540
rect 30318 232364 46318 240518
rect 57044 239300 58054 239500
rect 57044 238820 57198 239300
rect 57918 238820 58054 239300
rect 57044 238400 58054 238820
rect 60764 239300 61774 239500
rect 60764 238820 60918 239300
rect 61638 238820 61774 239300
rect 57064 232364 58032 238400
rect 60764 232528 61774 238820
rect 60730 232512 63776 232528
rect 73428 232512 89428 240376
rect 30318 231438 58072 232364
rect 30318 224318 46318 231438
rect 60730 231396 89428 232512
rect 73400 231288 89428 231396
rect 51806 228222 54366 229006
rect 51806 226544 52334 228222
rect 53754 226544 54366 228222
rect 51806 224276 54366 226544
rect 50782 208076 66782 224276
rect 73428 224176 89428 231288
rect 119442 232160 135442 240314
rect 146168 239096 147178 239296
rect 146168 238616 146322 239096
rect 147042 238616 147178 239096
rect 146168 238196 147178 238616
rect 149888 239096 150898 239296
rect 149888 238616 150042 239096
rect 150762 238616 150898 239096
rect 146188 232160 147156 238196
rect 149888 232324 150898 238616
rect 149854 232308 152900 232324
rect 162552 232308 178552 240172
rect 119442 231234 147196 232160
rect 119442 224114 135442 231234
rect 149854 231192 178552 232308
rect 162524 231084 178552 231192
rect 140930 228018 143490 228802
rect 140930 226340 141458 228018
rect 142878 226340 143490 228018
rect 140930 224072 143490 226340
rect 139906 207872 155906 224072
rect 162552 223972 178552 231084
rect 210696 231972 226696 240126
rect 237422 238908 238432 239108
rect 237422 238428 237576 238908
rect 238296 238428 238432 238908
rect 237422 238008 238432 238428
rect 241142 238908 242152 239108
rect 241142 238428 241296 238908
rect 242016 238428 242152 238908
rect 237442 231972 238410 238008
rect 241142 232136 242152 238428
rect 241108 232120 244154 232136
rect 253806 232120 269806 239984
rect 210696 231046 238450 231972
rect 210696 223926 226696 231046
rect 241108 231004 269806 232120
rect 253778 230896 269806 231004
rect 232184 227830 234744 228614
rect 232184 226152 232712 227830
rect 234132 226152 234744 227830
rect 232184 223884 234744 226152
rect 231160 207684 247160 223884
rect 253806 223784 269806 230896
rect 300318 232364 316318 240518
rect 327044 239300 328054 239500
rect 327044 238820 327198 239300
rect 327918 238820 328054 239300
rect 327044 238400 328054 238820
rect 330764 239300 331774 239500
rect 330764 238820 330918 239300
rect 331638 238820 331774 239300
rect 327064 232364 328032 238400
rect 330764 232528 331774 238820
rect 330730 232512 333776 232528
rect 343428 232512 359428 240376
rect 300318 231438 328072 232364
rect 300318 224318 316318 231438
rect 330730 231396 359428 232512
rect 343400 231288 359428 231396
rect 321806 228222 324366 229006
rect 321806 226544 322334 228222
rect 323754 226544 324366 228222
rect 321806 224276 324366 226544
rect 320782 208076 336782 224276
rect 343428 224176 359428 231288
rect 390318 232364 406318 240518
rect 417044 239300 418054 239500
rect 417044 238820 417198 239300
rect 417918 238820 418054 239300
rect 417044 238400 418054 238820
rect 420764 239300 421774 239500
rect 420764 238820 420918 239300
rect 421638 238820 421774 239300
rect 417064 232364 418032 238400
rect 420764 232528 421774 238820
rect 420730 232512 423776 232528
rect 433428 232512 449428 240376
rect 390318 231438 418072 232364
rect 390318 224318 406318 231438
rect 420730 231396 449428 232512
rect 433400 231288 449428 231396
rect 411806 228222 414366 229006
rect 411806 226544 412334 228222
rect 413754 226544 414366 228222
rect 411806 224276 414366 226544
rect 410782 208076 426782 224276
rect 433428 224176 449428 231288
rect 480318 232364 496318 240518
rect 507044 239300 508054 239500
rect 507044 238820 507198 239300
rect 507918 238820 508054 239300
rect 507044 238400 508054 238820
rect 510764 239300 511774 239500
rect 510764 238820 510918 239300
rect 511638 238820 511774 239300
rect 507064 232364 508032 238400
rect 510764 232528 511774 238820
rect 510730 232512 513776 232528
rect 523428 232512 539428 240376
rect 480318 231438 508072 232364
rect 480318 224318 496318 231438
rect 510730 231396 539428 232512
rect 523400 231288 539428 231396
rect 501806 228222 504366 229006
rect 501806 226544 502334 228222
rect 503754 226544 504366 228222
rect 501806 224276 504366 226544
rect 500782 208076 516782 224276
rect 523428 224176 539428 231288
rect 30332 166200 46332 171820
rect 30332 164940 58098 166200
rect 73518 166140 89518 171840
rect 72558 166124 89518 166140
rect 60790 165008 89518 166124
rect 60790 164992 63836 165008
rect 72558 165000 89518 165008
rect 30332 163040 46332 164940
rect 30198 162040 46338 163040
rect 30332 155620 46332 162040
rect 57124 159120 58092 164940
rect 57104 158700 58114 159120
rect 57104 158220 57258 158700
rect 57978 158220 58114 158700
rect 57104 158020 58114 158220
rect 60824 158700 61834 164992
rect 60824 158220 60978 158700
rect 61698 158220 61834 158700
rect 60824 158020 61834 158220
rect 73518 155640 89518 165000
rect 120332 166200 136332 171820
rect 120332 164940 148098 166200
rect 163518 166140 179518 171840
rect 162558 166124 179518 166140
rect 150790 165008 179518 166124
rect 150790 164992 153836 165008
rect 162558 165000 179518 165008
rect 120332 163040 136332 164940
rect 120198 162040 136338 163040
rect 120332 155620 136332 162040
rect 147124 159120 148092 164940
rect 147104 158700 148114 159120
rect 147104 158220 147258 158700
rect 147978 158220 148114 158700
rect 147104 158020 148114 158220
rect 150824 158700 151834 164992
rect 150824 158220 150978 158700
rect 151698 158220 151834 158700
rect 150824 158020 151834 158220
rect 163518 155640 179518 165000
rect 210332 166200 226332 171820
rect 210332 164940 238098 166200
rect 253518 166140 269518 171840
rect 252558 166124 269518 166140
rect 240790 165008 269518 166124
rect 240790 164992 243836 165008
rect 252558 165000 269518 165008
rect 210332 163040 226332 164940
rect 210198 162040 226338 163040
rect 210332 155620 226332 162040
rect 237124 159120 238092 164940
rect 237104 158700 238114 159120
rect 237104 158220 237258 158700
rect 237978 158220 238114 158700
rect 237104 158020 238114 158220
rect 240824 158700 241834 164992
rect 240824 158220 240978 158700
rect 241698 158220 241834 158700
rect 240824 158020 241834 158220
rect 253518 155640 269518 165000
rect 300332 166200 316332 171820
rect 300332 164940 328098 166200
rect 343518 166140 359518 171840
rect 342558 166124 359518 166140
rect 330790 165008 359518 166124
rect 330790 164992 333836 165008
rect 342558 165000 359518 165008
rect 300332 163040 316332 164940
rect 300198 162040 316338 163040
rect 300332 155620 316332 162040
rect 327124 159120 328092 164940
rect 327104 158700 328114 159120
rect 327104 158220 327258 158700
rect 327978 158220 328114 158700
rect 327104 158020 328114 158220
rect 330824 158700 331834 164992
rect 330824 158220 330978 158700
rect 331698 158220 331834 158700
rect 330824 158020 331834 158220
rect 343518 155640 359518 165000
rect 390332 166200 406332 171820
rect 390332 164940 418098 166200
rect 433518 166140 449518 171840
rect 432558 166124 449518 166140
rect 420790 165008 449518 166124
rect 420790 164992 423836 165008
rect 432558 165000 449518 165008
rect 390332 163040 406332 164940
rect 390198 162040 406338 163040
rect 390332 155620 406332 162040
rect 417124 159120 418092 164940
rect 417104 158700 418114 159120
rect 417104 158220 417258 158700
rect 417978 158220 418114 158700
rect 417104 158020 418114 158220
rect 420824 158700 421834 164992
rect 420824 158220 420978 158700
rect 421698 158220 421834 158700
rect 420824 158020 421834 158220
rect 433518 155640 449518 165000
rect 480332 166200 496332 171820
rect 480332 164940 508098 166200
rect 523518 166140 539518 171840
rect 522558 166124 539518 166140
rect 510790 165008 539518 166124
rect 510790 164992 513836 165008
rect 522558 165000 539518 165008
rect 480332 163040 496332 164940
rect 480198 162040 496338 163040
rect 480332 155620 496332 162040
rect 507124 159120 508092 164940
rect 507104 158700 508114 159120
rect 507104 158220 507258 158700
rect 507978 158220 508114 158700
rect 507104 158020 508114 158220
rect 510824 158700 511834 164992
rect 510824 158220 510978 158700
rect 511698 158220 511834 158700
rect 510824 158020 511834 158220
rect 523518 155640 539518 165000
rect 30398 145954 46398 153140
rect 73428 146094 89428 153106
rect 30398 145950 53488 145954
rect 30398 145260 53546 145950
rect 30398 144940 53194 145260
rect 53514 144940 53546 145260
rect 30398 144664 53546 144940
rect 66398 145724 89428 146094
rect 66398 145090 66566 145724
rect 67218 145090 89428 145724
rect 30398 136940 46398 144664
rect 66398 144554 89428 145090
rect 73428 136906 89428 144554
rect 120398 145954 136398 153140
rect 163428 146094 179428 153106
rect 120398 145950 143488 145954
rect 120398 145260 143546 145950
rect 120398 144940 143194 145260
rect 143514 144940 143546 145260
rect 120398 144664 143546 144940
rect 156398 145724 179428 146094
rect 156398 145090 156566 145724
rect 157218 145090 179428 145724
rect 120398 136940 136398 144664
rect 156398 144554 179428 145090
rect 163428 136906 179428 144554
rect 210398 145954 226398 153140
rect 253428 146094 269428 153106
rect 210398 145950 233488 145954
rect 210398 145260 233546 145950
rect 210398 144940 233194 145260
rect 233514 144940 233546 145260
rect 210398 144664 233546 144940
rect 246398 145724 269428 146094
rect 246398 145090 246566 145724
rect 247218 145090 269428 145724
rect 210398 136940 226398 144664
rect 246398 144554 269428 145090
rect 253428 136906 269428 144554
rect 300398 145954 316398 153140
rect 343428 146094 359428 153106
rect 300398 145950 323488 145954
rect 300398 145260 323546 145950
rect 300398 144940 323194 145260
rect 323514 144940 323546 145260
rect 300398 144664 323546 144940
rect 336398 145724 359428 146094
rect 336398 145090 336566 145724
rect 337218 145090 359428 145724
rect 300398 136940 316398 144664
rect 336398 144554 359428 145090
rect 343428 136906 359428 144554
rect 390398 145954 406398 153140
rect 433428 146094 449428 153106
rect 390398 145950 413488 145954
rect 390398 145260 413546 145950
rect 390398 144940 413194 145260
rect 413514 144940 413546 145260
rect 390398 144664 413546 144940
rect 426398 145724 449428 146094
rect 426398 145090 426566 145724
rect 427218 145090 449428 145724
rect 390398 136940 406398 144664
rect 426398 144554 449428 145090
rect 433428 136906 449428 144554
rect 480398 145954 496398 153140
rect 523428 146094 539428 153106
rect 480398 145950 503488 145954
rect 480398 145260 503546 145950
rect 480398 144940 503194 145260
rect 503514 144940 503546 145260
rect 480398 144664 503546 144940
rect 516398 145724 539428 146094
rect 516398 145090 516566 145724
rect 517218 145090 539428 145724
rect 480398 136940 496398 144664
rect 516398 144554 539428 145090
rect 523428 136906 539428 144554
rect 30318 126264 46318 134418
rect 57044 133200 58054 133400
rect 57044 132720 57198 133200
rect 57918 132720 58054 133200
rect 57044 132300 58054 132720
rect 60764 133200 61774 133400
rect 60764 132720 60918 133200
rect 61638 132720 61774 133200
rect 57064 126264 58032 132300
rect 60764 126428 61774 132720
rect 60730 126412 63776 126428
rect 73428 126412 89428 134276
rect 30318 125338 58072 126264
rect 30318 118218 46318 125338
rect 60730 125296 89428 126412
rect 73400 125188 89428 125296
rect 73428 118076 89428 125188
rect 120318 126264 136318 134418
rect 147044 133200 148054 133400
rect 147044 132720 147198 133200
rect 147918 132720 148054 133200
rect 147044 132300 148054 132720
rect 150764 133200 151774 133400
rect 150764 132720 150918 133200
rect 151638 132720 151774 133200
rect 147064 126264 148032 132300
rect 150764 126428 151774 132720
rect 150730 126412 153776 126428
rect 163428 126412 179428 134276
rect 120318 125338 148072 126264
rect 120318 118218 136318 125338
rect 150730 125296 179428 126412
rect 163400 125188 179428 125296
rect 163428 118076 179428 125188
rect 210318 126264 226318 134418
rect 237044 133200 238054 133400
rect 237044 132720 237198 133200
rect 237918 132720 238054 133200
rect 237044 132300 238054 132720
rect 240764 133200 241774 133400
rect 240764 132720 240918 133200
rect 241638 132720 241774 133200
rect 237064 126264 238032 132300
rect 240764 126428 241774 132720
rect 240730 126412 243776 126428
rect 253428 126412 269428 134276
rect 210318 125338 238072 126264
rect 210318 118218 226318 125338
rect 240730 125296 269428 126412
rect 253400 125188 269428 125296
rect 253428 118076 269428 125188
rect 300318 126264 316318 134418
rect 327044 133200 328054 133400
rect 327044 132720 327198 133200
rect 327918 132720 328054 133200
rect 327044 132300 328054 132720
rect 330764 133200 331774 133400
rect 330764 132720 330918 133200
rect 331638 132720 331774 133200
rect 327064 126264 328032 132300
rect 330764 126428 331774 132720
rect 330730 126412 333776 126428
rect 343428 126412 359428 134276
rect 300318 125338 328072 126264
rect 300318 118218 316318 125338
rect 330730 125296 359428 126412
rect 343400 125188 359428 125296
rect 343428 118076 359428 125188
rect 390318 126264 406318 134418
rect 417044 133200 418054 133400
rect 417044 132720 417198 133200
rect 417918 132720 418054 133200
rect 417044 132300 418054 132720
rect 420764 133200 421774 133400
rect 420764 132720 420918 133200
rect 421638 132720 421774 133200
rect 417064 126264 418032 132300
rect 420764 126428 421774 132720
rect 420730 126412 423776 126428
rect 433428 126412 449428 134276
rect 390318 125338 418072 126264
rect 390318 118218 406318 125338
rect 420730 125296 449428 126412
rect 433400 125188 449428 125296
rect 433428 118076 449428 125188
rect 480318 126264 496318 134418
rect 507044 133200 508054 133400
rect 507044 132720 507198 133200
rect 507918 132720 508054 133200
rect 507044 132300 508054 132720
rect 510764 133200 511774 133400
rect 510764 132720 510918 133200
rect 511638 132720 511774 133200
rect 507064 126264 508032 132300
rect 510764 126428 511774 132720
rect 510730 126412 513776 126428
rect 523428 126412 539428 134276
rect 480318 125338 508072 126264
rect 480318 118218 496318 125338
rect 510730 125296 539428 126412
rect 523400 125188 539428 125296
rect 523428 118076 539428 125188
rect 30332 76200 46332 81820
rect 30332 74940 58098 76200
rect 73518 76140 89518 81840
rect 72558 76124 89518 76140
rect 60790 75008 89518 76124
rect 60790 74992 63836 75008
rect 72558 75000 89518 75008
rect 30332 73040 46332 74940
rect 30198 72040 46338 73040
rect 30332 65620 46332 72040
rect 57124 69120 58092 74940
rect 57104 68700 58114 69120
rect 57104 68220 57258 68700
rect 57978 68220 58114 68700
rect 57104 68020 58114 68220
rect 60824 68700 61834 74992
rect 60824 68220 60978 68700
rect 61698 68220 61834 68700
rect 60824 68020 61834 68220
rect 73518 65640 89518 75000
rect 120332 76200 136332 81820
rect 120332 74940 148098 76200
rect 163518 76140 179518 81840
rect 162558 76124 179518 76140
rect 150790 75008 179518 76124
rect 150790 74992 153836 75008
rect 162558 75000 179518 75008
rect 120332 73040 136332 74940
rect 120198 72040 136338 73040
rect 120332 65620 136332 72040
rect 147124 69120 148092 74940
rect 147104 68700 148114 69120
rect 147104 68220 147258 68700
rect 147978 68220 148114 68700
rect 147104 68020 148114 68220
rect 150824 68700 151834 74992
rect 150824 68220 150978 68700
rect 151698 68220 151834 68700
rect 150824 68020 151834 68220
rect 163518 65640 179518 75000
rect 210332 76200 226332 81820
rect 210332 74940 238098 76200
rect 253518 76140 269518 81840
rect 252558 76124 269518 76140
rect 240790 75008 269518 76124
rect 240790 74992 243836 75008
rect 252558 75000 269518 75008
rect 210332 73040 226332 74940
rect 210198 72040 226338 73040
rect 210332 65620 226332 72040
rect 237124 69120 238092 74940
rect 237104 68700 238114 69120
rect 237104 68220 237258 68700
rect 237978 68220 238114 68700
rect 237104 68020 238114 68220
rect 240824 68700 241834 74992
rect 240824 68220 240978 68700
rect 241698 68220 241834 68700
rect 240824 68020 241834 68220
rect 253518 65640 269518 75000
rect 300332 76200 316332 81820
rect 300332 74940 328098 76200
rect 343518 76140 359518 81840
rect 342558 76124 359518 76140
rect 330790 75008 359518 76124
rect 330790 74992 333836 75008
rect 342558 75000 359518 75008
rect 300332 73040 316332 74940
rect 300198 72040 316338 73040
rect 300332 65620 316332 72040
rect 327124 69120 328092 74940
rect 327104 68700 328114 69120
rect 327104 68220 327258 68700
rect 327978 68220 328114 68700
rect 327104 68020 328114 68220
rect 330824 68700 331834 74992
rect 330824 68220 330978 68700
rect 331698 68220 331834 68700
rect 330824 68020 331834 68220
rect 343518 65640 359518 75000
rect 390332 76200 406332 81820
rect 390332 74940 418098 76200
rect 433518 76140 449518 81840
rect 432558 76124 449518 76140
rect 420790 75008 449518 76124
rect 420790 74992 423836 75008
rect 432558 75000 449518 75008
rect 390332 73040 406332 74940
rect 390198 72040 406338 73040
rect 390332 65620 406332 72040
rect 417124 69120 418092 74940
rect 417104 68700 418114 69120
rect 417104 68220 417258 68700
rect 417978 68220 418114 68700
rect 417104 68020 418114 68220
rect 420824 68700 421834 74992
rect 420824 68220 420978 68700
rect 421698 68220 421834 68700
rect 420824 68020 421834 68220
rect 433518 65640 449518 75000
rect 480332 76200 496332 81820
rect 480332 74940 508098 76200
rect 523518 76140 539518 81840
rect 522558 76124 539518 76140
rect 510790 75008 539518 76124
rect 510790 74992 513836 75008
rect 522558 75000 539518 75008
rect 480332 73040 496332 74940
rect 480198 72040 496338 73040
rect 480332 65620 496332 72040
rect 507124 69120 508092 74940
rect 507104 68700 508114 69120
rect 507104 68220 507258 68700
rect 507978 68220 508114 68700
rect 507104 68020 508114 68220
rect 510824 68700 511834 74992
rect 510824 68220 510978 68700
rect 511698 68220 511834 68700
rect 510824 68020 511834 68220
rect 523518 65640 539518 75000
rect 30398 55954 46398 63140
rect 73428 56094 89428 63106
rect 30398 55950 53488 55954
rect 30398 55260 53546 55950
rect 30398 54940 53194 55260
rect 53514 54940 53546 55260
rect 30398 54664 53546 54940
rect 66398 55724 89428 56094
rect 66398 55090 66566 55724
rect 67218 55090 89428 55724
rect 30398 46940 46398 54664
rect 66398 54554 89428 55090
rect 73428 46906 89428 54554
rect 120398 55954 136398 63140
rect 163428 56094 179428 63106
rect 120398 55950 143488 55954
rect 120398 55260 143546 55950
rect 120398 54940 143194 55260
rect 143514 54940 143546 55260
rect 120398 54664 143546 54940
rect 156398 55724 179428 56094
rect 156398 55090 156566 55724
rect 157218 55090 179428 55724
rect 120398 46940 136398 54664
rect 156398 54554 179428 55090
rect 163428 46906 179428 54554
rect 210398 55954 226398 63140
rect 253428 56094 269428 63106
rect 210398 55950 233488 55954
rect 210398 55260 233546 55950
rect 210398 54940 233194 55260
rect 233514 54940 233546 55260
rect 210398 54664 233546 54940
rect 246398 55724 269428 56094
rect 246398 55090 246566 55724
rect 247218 55090 269428 55724
rect 210398 46940 226398 54664
rect 246398 54554 269428 55090
rect 253428 46906 269428 54554
rect 300398 55954 316398 63140
rect 343428 56094 359428 63106
rect 300398 55950 323488 55954
rect 300398 55260 323546 55950
rect 300398 54940 323194 55260
rect 323514 54940 323546 55260
rect 300398 54664 323546 54940
rect 336398 55724 359428 56094
rect 336398 55090 336566 55724
rect 337218 55090 359428 55724
rect 300398 46940 316398 54664
rect 336398 54554 359428 55090
rect 343428 46906 359428 54554
rect 390398 55954 406398 63140
rect 433428 56094 449428 63106
rect 390398 55950 413488 55954
rect 390398 55260 413546 55950
rect 390398 54940 413194 55260
rect 413514 54940 413546 55260
rect 390398 54664 413546 54940
rect 426398 55724 449428 56094
rect 426398 55090 426566 55724
rect 427218 55090 449428 55724
rect 390398 46940 406398 54664
rect 426398 54554 449428 55090
rect 433428 46906 449428 54554
rect 480398 55954 496398 63140
rect 523428 56094 539428 63106
rect 480398 55950 503488 55954
rect 480398 55260 503546 55950
rect 480398 54940 503194 55260
rect 503514 54940 503546 55260
rect 480398 54664 503546 54940
rect 516398 55724 539428 56094
rect 516398 55090 516566 55724
rect 517218 55090 539428 55724
rect 480398 46940 496398 54664
rect 516398 54554 539428 55090
rect 523428 46906 539428 54554
rect 30318 36264 46318 44418
rect 57044 43200 58054 43400
rect 57044 42720 57198 43200
rect 57918 42720 58054 43200
rect 57044 42300 58054 42720
rect 60764 43200 61774 43400
rect 60764 42720 60918 43200
rect 61638 42720 61774 43200
rect 57064 36264 58032 42300
rect 60764 36428 61774 42720
rect 60730 36412 63776 36428
rect 73428 36412 89428 44276
rect 30318 35338 58072 36264
rect 30318 28218 46318 35338
rect 60730 35296 89428 36412
rect 73400 35188 89428 35296
rect 73428 28076 89428 35188
rect 120318 36264 136318 44418
rect 147044 43200 148054 43400
rect 147044 42720 147198 43200
rect 147918 42720 148054 43200
rect 147044 42300 148054 42720
rect 150764 43200 151774 43400
rect 150764 42720 150918 43200
rect 151638 42720 151774 43200
rect 147064 36264 148032 42300
rect 150764 36428 151774 42720
rect 150730 36412 153776 36428
rect 163428 36412 179428 44276
rect 120318 35338 148072 36264
rect 120318 28218 136318 35338
rect 150730 35296 179428 36412
rect 163400 35188 179428 35296
rect 163428 28076 179428 35188
rect 210318 36264 226318 44418
rect 237044 43200 238054 43400
rect 237044 42720 237198 43200
rect 237918 42720 238054 43200
rect 237044 42300 238054 42720
rect 240764 43200 241774 43400
rect 240764 42720 240918 43200
rect 241638 42720 241774 43200
rect 237064 36264 238032 42300
rect 240764 36428 241774 42720
rect 240730 36412 243776 36428
rect 253428 36412 269428 44276
rect 210318 35338 238072 36264
rect 210318 28218 226318 35338
rect 240730 35296 269428 36412
rect 253400 35188 269428 35296
rect 253428 28076 269428 35188
rect 300318 36264 316318 44418
rect 327044 43200 328054 43400
rect 327044 42720 327198 43200
rect 327918 42720 328054 43200
rect 327044 42300 328054 42720
rect 330764 43200 331774 43400
rect 330764 42720 330918 43200
rect 331638 42720 331774 43200
rect 327064 36264 328032 42300
rect 330764 36428 331774 42720
rect 330730 36412 333776 36428
rect 343428 36412 359428 44276
rect 300318 35338 328072 36264
rect 300318 28218 316318 35338
rect 330730 35296 359428 36412
rect 343400 35188 359428 35296
rect 343428 28076 359428 35188
rect 390318 36264 406318 44418
rect 417044 43200 418054 43400
rect 417044 42720 417198 43200
rect 417918 42720 418054 43200
rect 417044 42300 418054 42720
rect 420764 43200 421774 43400
rect 420764 42720 420918 43200
rect 421638 42720 421774 43200
rect 417064 36264 418032 42300
rect 420764 36428 421774 42720
rect 420730 36412 423776 36428
rect 433428 36412 449428 44276
rect 390318 35338 418072 36264
rect 390318 28218 406318 35338
rect 420730 35296 449428 36412
rect 433400 35188 449428 35296
rect 433428 28076 449428 35188
rect 480318 36264 496318 44418
rect 507044 43200 508054 43400
rect 507044 42720 507198 43200
rect 507918 42720 508054 43200
rect 507044 42300 508054 42720
rect 510764 43200 511774 43400
rect 510764 42720 510918 43200
rect 511638 42720 511774 43200
rect 507064 36264 508032 42300
rect 510764 36428 511774 42720
rect 510730 36412 513776 36428
rect 523428 36412 539428 44276
rect 480318 35338 508072 36264
rect 480318 28218 496318 35338
rect 510730 35296 539428 36412
rect 523400 35188 539428 35296
rect 523428 28076 539428 35188
<< glass >>
rect 30798 665840 45932 681420
rect 73918 666040 88998 681440
rect 120798 665840 135932 681420
rect 163918 666040 178998 681440
rect 210798 665840 225932 681420
rect 253918 666040 268998 681440
rect 300600 667764 315734 683344
rect 343720 667964 358800 683364
rect 390600 667764 405734 683344
rect 433720 667964 448800 683364
rect 480600 667764 495734 683344
rect 523720 667964 538800 683364
rect 30798 647340 45998 662740
rect 73828 647306 89028 662706
rect 120798 647340 135998 662740
rect 163828 647306 179028 662706
rect 210798 647340 225998 662740
rect 253828 647306 269028 662706
rect 300600 649264 315800 664664
rect 343630 649230 358830 664630
rect 390600 649264 405800 664664
rect 433630 649230 448830 664630
rect 480600 649264 495800 664664
rect 523630 649230 538830 664630
rect 30718 628640 45918 644020
rect 73828 628476 89028 643876
rect 120718 628640 135918 644020
rect 163828 628476 179028 643876
rect 210718 628640 225918 644020
rect 253828 628476 269028 643876
rect 300520 630564 315720 645944
rect 343630 630400 358830 645800
rect 390520 630564 405720 645944
rect 433630 630400 448830 645800
rect 480520 630564 495720 645944
rect 523630 630400 538830 645800
rect 30798 590840 45932 606420
rect 73918 591040 88998 606440
rect 120798 590840 135932 606420
rect 163918 591040 178998 606440
rect 210798 590840 225932 606420
rect 253918 591040 268998 606440
rect 300798 590840 315932 606420
rect 343918 591040 358998 606440
rect 390600 592764 405734 608344
rect 433720 592964 448800 608364
rect 480600 592764 495734 608344
rect 523720 592964 538800 608364
rect 30798 572340 45998 587740
rect 73828 572306 89028 587706
rect 120798 572340 135998 587740
rect 163828 572306 179028 587706
rect 210798 572340 225998 587740
rect 253828 572306 269028 587706
rect 300798 572340 315998 587740
rect 343828 572306 359028 587706
rect 390600 574264 405800 589664
rect 433630 574230 448830 589630
rect 480600 574264 495800 589664
rect 523630 574230 538830 589630
rect 30718 553640 45918 569020
rect 73828 553476 89028 568876
rect 120718 553640 135918 569020
rect 163828 553476 179028 568876
rect 210718 553640 225918 569020
rect 253828 553476 269028 568876
rect 300718 553640 315918 569020
rect 343828 553476 359028 568876
rect 390520 555564 405720 570944
rect 433630 555400 448830 570800
rect 480520 555564 495720 570944
rect 523630 555400 538830 570800
rect 51598 518340 66998 533740
rect 141598 518340 156998 533740
rect 231598 518340 246998 533740
rect 321598 518340 336998 533740
rect 411598 518340 426998 533740
rect 501598 518340 516998 533740
rect 30798 501940 45932 517520
rect 73918 502140 88998 517540
rect 120798 501940 135932 517520
rect 163918 502140 178998 517540
rect 210798 501940 225932 517520
rect 253918 502140 268998 517540
rect 300798 501940 315932 517520
rect 343918 502140 358998 517540
rect 390798 501940 405932 517520
rect 433918 502140 448998 517540
rect 480798 501940 495932 517520
rect 523918 502140 538998 517540
rect 30798 483440 45998 498840
rect 73828 483406 89028 498806
rect 120798 483440 135998 498840
rect 163828 483406 179028 498806
rect 210798 483440 225998 498840
rect 253828 483406 269028 498806
rect 300798 483440 315998 498840
rect 343828 483406 359028 498806
rect 390798 483440 405998 498840
rect 433828 483406 449028 498806
rect 480798 483440 495998 498840
rect 523828 483406 539028 498806
rect 30718 464740 45918 480120
rect 73828 464576 89028 479976
rect 120718 464740 135918 480120
rect 163828 464576 179028 479976
rect 210718 464740 225918 480120
rect 253828 464576 269028 479976
rect 300718 464740 315918 480120
rect 343828 464576 359028 479976
rect 390718 464740 405918 480120
rect 433828 464576 449028 479976
rect 480718 464740 495918 480120
rect 523828 464576 539028 479976
rect 51198 448340 66398 463940
rect 141198 448340 156398 463940
rect 231198 448340 246398 463940
rect 321198 448340 336398 463940
rect 411198 448340 426398 463940
rect 501198 448340 516398 463940
rect 51598 398340 66998 413740
rect 141598 398340 156998 413740
rect 231598 398340 246998 413740
rect 321598 398340 336998 413740
rect 411598 398340 426998 413740
rect 501598 398340 516998 413740
rect 30798 381940 45932 397520
rect 73918 382140 88998 397540
rect 120798 381940 135932 397520
rect 163918 382140 178998 397540
rect 210798 381940 225932 397520
rect 253918 382140 268998 397540
rect 300798 381940 315932 397520
rect 343918 382140 358998 397540
rect 390798 381940 405932 397520
rect 433918 382140 448998 397540
rect 480798 381940 495932 397520
rect 523918 382140 538998 397540
rect 30798 363440 45998 378840
rect 73828 363406 89028 378806
rect 120798 363440 135998 378840
rect 163828 363406 179028 378806
rect 210798 363440 225998 378840
rect 253828 363406 269028 378806
rect 300798 363440 315998 378840
rect 343828 363406 359028 378806
rect 390798 363440 405998 378840
rect 433828 363406 449028 378806
rect 480798 363440 495998 378840
rect 523828 363406 539028 378806
rect 30718 344740 45918 360120
rect 73828 344576 89028 359976
rect 120718 344740 135918 360120
rect 163828 344576 179028 359976
rect 210718 344740 225918 360120
rect 253828 344576 269028 359976
rect 300718 344740 315918 360120
rect 343828 344576 359028 359976
rect 390718 344740 405918 360120
rect 433828 344576 449028 359976
rect 480718 344740 495918 360120
rect 523828 344576 539028 359976
rect 51198 328340 66398 343940
rect 141198 328340 156398 343940
rect 231198 328340 246398 343940
rect 321198 328340 336398 343940
rect 411198 328340 426398 343940
rect 501198 328340 516398 343940
rect 51598 278340 66998 293740
rect 140722 278136 156122 293536
rect 231976 277948 247376 293348
rect 321598 278340 336998 293740
rect 411598 278340 426998 293740
rect 501598 278340 516998 293740
rect 30798 261940 45932 277520
rect 73918 262140 88998 277540
rect 119922 261736 135056 277316
rect 163042 261936 178122 277336
rect 211176 261548 226310 277128
rect 254296 261748 269376 277148
rect 300798 261940 315932 277520
rect 343918 262140 358998 277540
rect 390798 261940 405932 277520
rect 433918 262140 448998 277540
rect 480798 261940 495932 277520
rect 523918 262140 538998 277540
rect 30798 243440 45998 258840
rect 73828 243406 89028 258806
rect 119922 243236 135122 258636
rect 162952 243202 178152 258602
rect 211176 243048 226376 258448
rect 254206 243014 269406 258414
rect 300798 243440 315998 258840
rect 343828 243406 359028 258806
rect 390798 243440 405998 258840
rect 433828 243406 449028 258806
rect 480798 243440 495998 258840
rect 523828 243406 539028 258806
rect 30718 224740 45918 240120
rect 73828 224576 89028 239976
rect 119842 224536 135042 239916
rect 162952 224372 178152 239772
rect 211096 224348 226296 239728
rect 254206 224184 269406 239584
rect 300718 224740 315918 240120
rect 343828 224576 359028 239976
rect 390718 224740 405918 240120
rect 433828 224576 449028 239976
rect 480718 224740 495918 240120
rect 523828 224576 539028 239976
rect 51198 208340 66398 223940
rect 140322 208136 155522 223736
rect 231576 207948 246776 223548
rect 321198 208340 336398 223940
rect 411198 208340 426398 223940
rect 501198 208340 516398 223940
rect 30798 155840 45932 171420
rect 73918 156040 88998 171440
rect 120798 155840 135932 171420
rect 163918 156040 178998 171440
rect 210798 155840 225932 171420
rect 253918 156040 268998 171440
rect 300798 155840 315932 171420
rect 343918 156040 358998 171440
rect 390798 155840 405932 171420
rect 433918 156040 448998 171440
rect 480798 155840 495932 171420
rect 523918 156040 538998 171440
rect 30798 137340 45998 152740
rect 73828 137306 89028 152706
rect 120798 137340 135998 152740
rect 163828 137306 179028 152706
rect 210798 137340 225998 152740
rect 253828 137306 269028 152706
rect 300798 137340 315998 152740
rect 343828 137306 359028 152706
rect 390798 137340 405998 152740
rect 433828 137306 449028 152706
rect 480798 137340 495998 152740
rect 523828 137306 539028 152706
rect 30718 118640 45918 134020
rect 73828 118476 89028 133876
rect 120718 118640 135918 134020
rect 163828 118476 179028 133876
rect 210718 118640 225918 134020
rect 253828 118476 269028 133876
rect 300718 118640 315918 134020
rect 343828 118476 359028 133876
rect 390718 118640 405918 134020
rect 433828 118476 449028 133876
rect 480718 118640 495918 134020
rect 523828 118476 539028 133876
rect 30798 65840 45932 81420
rect 73918 66040 88998 81440
rect 120798 65840 135932 81420
rect 163918 66040 178998 81440
rect 210798 65840 225932 81420
rect 253918 66040 268998 81440
rect 300798 65840 315932 81420
rect 343918 66040 358998 81440
rect 390798 65840 405932 81420
rect 433918 66040 448998 81440
rect 480798 65840 495932 81420
rect 523918 66040 538998 81440
rect 30798 47340 45998 62740
rect 73828 47306 89028 62706
rect 120798 47340 135998 62740
rect 163828 47306 179028 62706
rect 210798 47340 225998 62740
rect 253828 47306 269028 62706
rect 300798 47340 315998 62740
rect 343828 47306 359028 62706
rect 390798 47340 405998 62740
rect 433828 47306 449028 62706
rect 480798 47340 495998 62740
rect 523828 47306 539028 62706
rect 30718 28640 45918 44020
rect 73828 28476 89028 43876
rect 120718 28640 135918 44020
rect 163828 28476 179028 43876
rect 210718 28640 225918 44020
rect 253828 28476 269028 43876
rect 300718 28640 315918 44020
rect 343828 28476 359028 43876
rect 390718 28640 405918 44020
rect 433828 28476 449028 43876
rect 480718 28640 495918 44020
rect 523828 28476 539028 43876
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1400 0 0 0 gpio_analog[0]
port 1 nsew
flabel metal3 s -800 381864 480 381976 0 FreeSans 1400 0 0 0 gpio_analog[10]
port 2 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 1400 0 0 0 gpio_analog[11]
port 3 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1400 0 0 0 gpio_analog[12]
port 4 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 1400 0 0 0 gpio_analog[13]
port 5 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 1400 0 0 0 gpio_analog[14]
port 6 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 1400 0 0 0 gpio_analog[15]
port 7 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 1400 0 0 0 gpio_analog[16]
port 8 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 1400 0 0 0 gpio_analog[17]
port 9 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1400 0 0 0 gpio_analog[1]
port 10 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1400 0 0 0 gpio_analog[2]
port 11 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1400 0 0 0 gpio_analog[3]
port 12 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1400 0 0 0 gpio_analog[4]
port 13 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1400 0 0 0 gpio_analog[5]
port 14 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1400 0 0 0 gpio_analog[6]
port 15 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 1400 0 0 0 gpio_analog[7]
port 16 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 1400 0 0 0 gpio_analog[8]
port 17 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 1400 0 0 0 gpio_analog[9]
port 18 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1400 0 0 0 gpio_noesd[0]
port 19 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 1400 0 0 0 gpio_noesd[10]
port 20 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 1400 0 0 0 gpio_noesd[11]
port 21 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1400 0 0 0 gpio_noesd[12]
port 22 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 1400 0 0 0 gpio_noesd[13]
port 23 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 1400 0 0 0 gpio_noesd[14]
port 24 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 1400 0 0 0 gpio_noesd[15]
port 25 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 1400 0 0 0 gpio_noesd[16]
port 26 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 1400 0 0 0 gpio_noesd[17]
port 27 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1400 0 0 0 gpio_noesd[1]
port 28 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1400 0 0 0 gpio_noesd[2]
port 29 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1400 0 0 0 gpio_noesd[3]
port 30 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1400 0 0 0 gpio_noesd[4]
port 31 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1400 0 0 0 gpio_noesd[5]
port 32 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1400 0 0 0 gpio_noesd[6]
port 33 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 1400 0 0 0 gpio_noesd[7]
port 34 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 1400 0 0 0 gpio_noesd[8]
port 35 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 1400 0 0 0 gpio_noesd[9]
port 36 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1400 0 0 0 io_analog[0]
port 37 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1400 0 0 0 io_analog[10]
port 38 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 2400 180 0 0 io_analog[1]
port 39 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 2400 180 0 0 io_analog[2]
port 40 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 2400 180 0 0 io_analog[3]
port 41 nsew
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 2400 180 0 0 io_analog[7]
port 45 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 2400 180 0 0 io_analog[8]
port 46 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 2400 180 0 0 io_analog[9]
port 47 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 2400 180 0 0 io_clamp_high[0]
port 48 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 2400 180 0 0 io_clamp_high[1]
port 49 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 2400 180 0 0 io_clamp_high[2]
port 50 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 2400 180 0 0 io_clamp_low[0]
port 51 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 2400 180 0 0 io_clamp_low[1]
port 52 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 2400 180 0 0 io_clamp_low[2]
port 53 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1400 0 0 0 io_in[0]
port 54 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1400 0 0 0 io_in[10]
port 55 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1400 0 0 0 io_in[11]
port 56 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1400 0 0 0 io_in[12]
port 57 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1400 0 0 0 io_in[13]
port 58 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1400 0 0 0 io_in[14]
port 59 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 1400 0 0 0 io_in[15]
port 60 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1400 0 0 0 io_in[16]
port 61 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1400 0 0 0 io_in[17]
port 62 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1400 0 0 0 io_in[18]
port 63 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 1400 0 0 0 io_in[19]
port 64 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1400 0 0 0 io_in[1]
port 65 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 1400 0 0 0 io_in[20]
port 66 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 1400 0 0 0 io_in[21]
port 67 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 1400 0 0 0 io_in[22]
port 68 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 1400 0 0 0 io_in[23]
port 69 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 1400 0 0 0 io_in[24]
port 70 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 1400 0 0 0 io_in[25]
port 71 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 1400 0 0 0 io_in[26]
port 72 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1400 0 0 0 io_in[2]
port 73 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1400 0 0 0 io_in[3]
port 74 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1400 0 0 0 io_in[4]
port 75 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1400 0 0 0 io_in[5]
port 76 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1400 0 0 0 io_in[6]
port 77 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1400 0 0 0 io_in[7]
port 78 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1400 0 0 0 io_in[8]
port 79 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1400 0 0 0 io_in[9]
port 80 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1400 0 0 0 io_in_3v3[0]
port 81 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1400 0 0 0 io_in_3v3[10]
port 82 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1400 0 0 0 io_in_3v3[11]
port 83 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1400 0 0 0 io_in_3v3[12]
port 84 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1400 0 0 0 io_in_3v3[13]
port 85 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 1400 0 0 0 io_in_3v3[14]
port 86 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1400 0 0 0 io_in_3v3[15]
port 87 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 1400 0 0 0 io_in_3v3[16]
port 88 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 1400 0 0 0 io_in_3v3[17]
port 89 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 1400 0 0 0 io_in_3v3[18]
port 90 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 1400 0 0 0 io_in_3v3[19]
port 91 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1400 0 0 0 io_in_3v3[1]
port 92 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 1400 0 0 0 io_in_3v3[20]
port 93 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 1400 0 0 0 io_in_3v3[21]
port 94 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 1400 0 0 0 io_in_3v3[22]
port 95 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 1400 0 0 0 io_in_3v3[23]
port 96 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 1400 0 0 0 io_in_3v3[24]
port 97 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 1400 0 0 0 io_in_3v3[25]
port 98 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 1400 0 0 0 io_in_3v3[26]
port 99 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1400 0 0 0 io_in_3v3[2]
port 100 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1400 0 0 0 io_in_3v3[3]
port 101 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1400 0 0 0 io_in_3v3[4]
port 102 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1400 0 0 0 io_in_3v3[5]
port 103 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1400 0 0 0 io_in_3v3[6]
port 104 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1400 0 0 0 io_in_3v3[7]
port 105 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1400 0 0 0 io_in_3v3[8]
port 106 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1400 0 0 0 io_in_3v3[9]
port 107 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1400 0 0 0 io_oeb[0]
port 108 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1400 0 0 0 io_oeb[10]
port 109 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1400 0 0 0 io_oeb[11]
port 110 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1400 0 0 0 io_oeb[12]
port 111 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1400 0 0 0 io_oeb[13]
port 112 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 1400 0 0 0 io_oeb[14]
port 113 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 1400 0 0 0 io_oeb[15]
port 114 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 1400 0 0 0 io_oeb[16]
port 115 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 1400 0 0 0 io_oeb[17]
port 116 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 1400 0 0 0 io_oeb[18]
port 117 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 1400 0 0 0 io_oeb[19]
port 118 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1400 0 0 0 io_oeb[1]
port 119 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 1400 0 0 0 io_oeb[20]
port 120 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 1400 0 0 0 io_oeb[21]
port 121 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 1400 0 0 0 io_oeb[22]
port 122 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 1400 0 0 0 io_oeb[23]
port 123 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 1400 0 0 0 io_oeb[24]
port 124 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 1400 0 0 0 io_oeb[25]
port 125 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 1400 0 0 0 io_oeb[26]
port 126 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1400 0 0 0 io_oeb[2]
port 127 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1400 0 0 0 io_oeb[3]
port 128 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1400 0 0 0 io_oeb[4]
port 129 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1400 0 0 0 io_oeb[5]
port 130 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1400 0 0 0 io_oeb[6]
port 131 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1400 0 0 0 io_oeb[7]
port 132 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1400 0 0 0 io_oeb[8]
port 133 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1400 0 0 0 io_oeb[9]
port 134 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1400 0 0 0 io_out[0]
port 135 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1400 0 0 0 io_out[10]
port 136 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1400 0 0 0 io_out[11]
port 137 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1400 0 0 0 io_out[12]
port 138 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1400 0 0 0 io_out[13]
port 139 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 1400 0 0 0 io_out[14]
port 140 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 1400 0 0 0 io_out[15]
port 141 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 1400 0 0 0 io_out[16]
port 142 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 1400 0 0 0 io_out[17]
port 143 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 1400 0 0 0 io_out[18]
port 144 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 1400 0 0 0 io_out[19]
port 145 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1400 0 0 0 io_out[1]
port 146 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 1400 0 0 0 io_out[20]
port 147 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 1400 0 0 0 io_out[21]
port 148 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 1400 0 0 0 io_out[22]
port 149 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 1400 0 0 0 io_out[23]
port 150 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 1400 0 0 0 io_out[24]
port 151 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 1400 0 0 0 io_out[25]
port 152 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 1400 0 0 0 io_out[26]
port 153 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1400 0 0 0 io_out[2]
port 154 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1400 0 0 0 io_out[3]
port 155 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1400 0 0 0 io_out[4]
port 156 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1400 0 0 0 io_out[5]
port 157 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1400 0 0 0 io_out[6]
port 158 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1400 0 0 0 io_out[7]
port 159 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1400 0 0 0 io_out[8]
port 160 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1400 0 0 0 io_out[9]
port 161 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1400 90 0 0 la_data_in[0]
port 162 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1400 90 0 0 la_data_in[100]
port 163 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1400 90 0 0 la_data_in[101]
port 164 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1400 90 0 0 la_data_in[102]
port 165 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1400 90 0 0 la_data_in[103]
port 166 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1400 90 0 0 la_data_in[104]
port 167 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1400 90 0 0 la_data_in[105]
port 168 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1400 90 0 0 la_data_in[106]
port 169 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1400 90 0 0 la_data_in[107]
port 170 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1400 90 0 0 la_data_in[108]
port 171 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1400 90 0 0 la_data_in[109]
port 172 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1400 90 0 0 la_data_in[10]
port 173 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1400 90 0 0 la_data_in[110]
port 174 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1400 90 0 0 la_data_in[111]
port 175 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1400 90 0 0 la_data_in[112]
port 176 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1400 90 0 0 la_data_in[113]
port 177 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1400 90 0 0 la_data_in[114]
port 178 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1400 90 0 0 la_data_in[115]
port 179 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1400 90 0 0 la_data_in[116]
port 180 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1400 90 0 0 la_data_in[117]
port 181 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1400 90 0 0 la_data_in[118]
port 182 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1400 90 0 0 la_data_in[119]
port 183 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1400 90 0 0 la_data_in[11]
port 184 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1400 90 0 0 la_data_in[120]
port 185 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1400 90 0 0 la_data_in[121]
port 186 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1400 90 0 0 la_data_in[122]
port 187 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1400 90 0 0 la_data_in[123]
port 188 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1400 90 0 0 la_data_in[124]
port 189 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1400 90 0 0 la_data_in[125]
port 190 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1400 90 0 0 la_data_in[126]
port 191 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1400 90 0 0 la_data_in[127]
port 192 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1400 90 0 0 la_data_in[12]
port 193 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1400 90 0 0 la_data_in[13]
port 194 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1400 90 0 0 la_data_in[14]
port 195 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1400 90 0 0 la_data_in[15]
port 196 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1400 90 0 0 la_data_in[16]
port 197 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1400 90 0 0 la_data_in[17]
port 198 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1400 90 0 0 la_data_in[18]
port 199 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1400 90 0 0 la_data_in[19]
port 200 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1400 90 0 0 la_data_in[1]
port 201 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1400 90 0 0 la_data_in[20]
port 202 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1400 90 0 0 la_data_in[21]
port 203 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1400 90 0 0 la_data_in[22]
port 204 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1400 90 0 0 la_data_in[23]
port 205 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1400 90 0 0 la_data_in[24]
port 206 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1400 90 0 0 la_data_in[25]
port 207 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1400 90 0 0 la_data_in[26]
port 208 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1400 90 0 0 la_data_in[27]
port 209 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1400 90 0 0 la_data_in[28]
port 210 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1400 90 0 0 la_data_in[29]
port 211 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1400 90 0 0 la_data_in[2]
port 212 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1400 90 0 0 la_data_in[30]
port 213 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1400 90 0 0 la_data_in[31]
port 214 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1400 90 0 0 la_data_in[32]
port 215 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1400 90 0 0 la_data_in[33]
port 216 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1400 90 0 0 la_data_in[34]
port 217 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1400 90 0 0 la_data_in[35]
port 218 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1400 90 0 0 la_data_in[36]
port 219 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1400 90 0 0 la_data_in[37]
port 220 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1400 90 0 0 la_data_in[38]
port 221 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1400 90 0 0 la_data_in[39]
port 222 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1400 90 0 0 la_data_in[3]
port 223 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1400 90 0 0 la_data_in[40]
port 224 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1400 90 0 0 la_data_in[41]
port 225 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1400 90 0 0 la_data_in[42]
port 226 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1400 90 0 0 la_data_in[43]
port 227 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1400 90 0 0 la_data_in[44]
port 228 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1400 90 0 0 la_data_in[45]
port 229 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1400 90 0 0 la_data_in[46]
port 230 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1400 90 0 0 la_data_in[47]
port 231 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1400 90 0 0 la_data_in[48]
port 232 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1400 90 0 0 la_data_in[49]
port 233 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1400 90 0 0 la_data_in[4]
port 234 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1400 90 0 0 la_data_in[50]
port 235 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1400 90 0 0 la_data_in[51]
port 236 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1400 90 0 0 la_data_in[52]
port 237 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1400 90 0 0 la_data_in[53]
port 238 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1400 90 0 0 la_data_in[54]
port 239 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1400 90 0 0 la_data_in[55]
port 240 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1400 90 0 0 la_data_in[56]
port 241 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1400 90 0 0 la_data_in[57]
port 242 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1400 90 0 0 la_data_in[58]
port 243 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1400 90 0 0 la_data_in[59]
port 244 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1400 90 0 0 la_data_in[5]
port 245 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1400 90 0 0 la_data_in[60]
port 246 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1400 90 0 0 la_data_in[61]
port 247 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1400 90 0 0 la_data_in[62]
port 248 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1400 90 0 0 la_data_in[63]
port 249 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1400 90 0 0 la_data_in[64]
port 250 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1400 90 0 0 la_data_in[65]
port 251 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1400 90 0 0 la_data_in[66]
port 252 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1400 90 0 0 la_data_in[67]
port 253 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1400 90 0 0 la_data_in[68]
port 254 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1400 90 0 0 la_data_in[69]
port 255 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1400 90 0 0 la_data_in[6]
port 256 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1400 90 0 0 la_data_in[70]
port 257 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1400 90 0 0 la_data_in[71]
port 258 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1400 90 0 0 la_data_in[72]
port 259 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1400 90 0 0 la_data_in[73]
port 260 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1400 90 0 0 la_data_in[74]
port 261 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1400 90 0 0 la_data_in[75]
port 262 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1400 90 0 0 la_data_in[76]
port 263 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1400 90 0 0 la_data_in[77]
port 264 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1400 90 0 0 la_data_in[78]
port 265 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1400 90 0 0 la_data_in[79]
port 266 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1400 90 0 0 la_data_in[7]
port 267 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1400 90 0 0 la_data_in[80]
port 268 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1400 90 0 0 la_data_in[81]
port 269 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1400 90 0 0 la_data_in[82]
port 270 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1400 90 0 0 la_data_in[83]
port 271 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1400 90 0 0 la_data_in[84]
port 272 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1400 90 0 0 la_data_in[85]
port 273 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1400 90 0 0 la_data_in[86]
port 274 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1400 90 0 0 la_data_in[87]
port 275 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1400 90 0 0 la_data_in[88]
port 276 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1400 90 0 0 la_data_in[89]
port 277 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1400 90 0 0 la_data_in[8]
port 278 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1400 90 0 0 la_data_in[90]
port 279 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1400 90 0 0 la_data_in[91]
port 280 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1400 90 0 0 la_data_in[92]
port 281 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1400 90 0 0 la_data_in[93]
port 282 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1400 90 0 0 la_data_in[94]
port 283 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1400 90 0 0 la_data_in[95]
port 284 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1400 90 0 0 la_data_in[96]
port 285 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1400 90 0 0 la_data_in[97]
port 286 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1400 90 0 0 la_data_in[98]
port 287 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1400 90 0 0 la_data_in[99]
port 288 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1400 90 0 0 la_data_in[9]
port 289 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1400 90 0 0 la_data_out[0]
port 290 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1400 90 0 0 la_data_out[100]
port 291 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1400 90 0 0 la_data_out[101]
port 292 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1400 90 0 0 la_data_out[102]
port 293 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1400 90 0 0 la_data_out[103]
port 294 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1400 90 0 0 la_data_out[104]
port 295 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1400 90 0 0 la_data_out[105]
port 296 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1400 90 0 0 la_data_out[106]
port 297 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1400 90 0 0 la_data_out[107]
port 298 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1400 90 0 0 la_data_out[108]
port 299 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1400 90 0 0 la_data_out[109]
port 300 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1400 90 0 0 la_data_out[10]
port 301 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1400 90 0 0 la_data_out[110]
port 302 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1400 90 0 0 la_data_out[111]
port 303 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1400 90 0 0 la_data_out[112]
port 304 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1400 90 0 0 la_data_out[113]
port 305 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1400 90 0 0 la_data_out[114]
port 306 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1400 90 0 0 la_data_out[115]
port 307 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1400 90 0 0 la_data_out[116]
port 308 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1400 90 0 0 la_data_out[117]
port 309 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1400 90 0 0 la_data_out[118]
port 310 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1400 90 0 0 la_data_out[119]
port 311 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1400 90 0 0 la_data_out[11]
port 312 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1400 90 0 0 la_data_out[120]
port 313 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1400 90 0 0 la_data_out[121]
port 314 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1400 90 0 0 la_data_out[122]
port 315 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1400 90 0 0 la_data_out[123]
port 316 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1400 90 0 0 la_data_out[124]
port 317 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1400 90 0 0 la_data_out[125]
port 318 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1400 90 0 0 la_data_out[126]
port 319 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1400 90 0 0 la_data_out[127]
port 320 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1400 90 0 0 la_data_out[12]
port 321 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1400 90 0 0 la_data_out[13]
port 322 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1400 90 0 0 la_data_out[14]
port 323 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1400 90 0 0 la_data_out[15]
port 324 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1400 90 0 0 la_data_out[16]
port 325 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1400 90 0 0 la_data_out[17]
port 326 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1400 90 0 0 la_data_out[18]
port 327 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1400 90 0 0 la_data_out[19]
port 328 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1400 90 0 0 la_data_out[1]
port 329 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1400 90 0 0 la_data_out[20]
port 330 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1400 90 0 0 la_data_out[21]
port 331 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1400 90 0 0 la_data_out[22]
port 332 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1400 90 0 0 la_data_out[23]
port 333 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1400 90 0 0 la_data_out[24]
port 334 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1400 90 0 0 la_data_out[25]
port 335 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1400 90 0 0 la_data_out[26]
port 336 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1400 90 0 0 la_data_out[27]
port 337 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1400 90 0 0 la_data_out[28]
port 338 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1400 90 0 0 la_data_out[29]
port 339 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1400 90 0 0 la_data_out[2]
port 340 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1400 90 0 0 la_data_out[30]
port 341 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1400 90 0 0 la_data_out[31]
port 342 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1400 90 0 0 la_data_out[32]
port 343 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1400 90 0 0 la_data_out[33]
port 344 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1400 90 0 0 la_data_out[34]
port 345 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1400 90 0 0 la_data_out[35]
port 346 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1400 90 0 0 la_data_out[36]
port 347 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1400 90 0 0 la_data_out[37]
port 348 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1400 90 0 0 la_data_out[38]
port 349 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1400 90 0 0 la_data_out[39]
port 350 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1400 90 0 0 la_data_out[3]
port 351 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1400 90 0 0 la_data_out[40]
port 352 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1400 90 0 0 la_data_out[41]
port 353 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1400 90 0 0 la_data_out[42]
port 354 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1400 90 0 0 la_data_out[43]
port 355 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1400 90 0 0 la_data_out[44]
port 356 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1400 90 0 0 la_data_out[45]
port 357 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1400 90 0 0 la_data_out[46]
port 358 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1400 90 0 0 la_data_out[47]
port 359 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1400 90 0 0 la_data_out[48]
port 360 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1400 90 0 0 la_data_out[49]
port 361 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1400 90 0 0 la_data_out[4]
port 362 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1400 90 0 0 la_data_out[50]
port 363 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1400 90 0 0 la_data_out[51]
port 364 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1400 90 0 0 la_data_out[52]
port 365 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1400 90 0 0 la_data_out[53]
port 366 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1400 90 0 0 la_data_out[54]
port 367 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1400 90 0 0 la_data_out[55]
port 368 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1400 90 0 0 la_data_out[56]
port 369 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1400 90 0 0 la_data_out[57]
port 370 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1400 90 0 0 la_data_out[58]
port 371 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1400 90 0 0 la_data_out[59]
port 372 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1400 90 0 0 la_data_out[5]
port 373 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1400 90 0 0 la_data_out[60]
port 374 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1400 90 0 0 la_data_out[61]
port 375 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1400 90 0 0 la_data_out[62]
port 376 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1400 90 0 0 la_data_out[63]
port 377 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1400 90 0 0 la_data_out[64]
port 378 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1400 90 0 0 la_data_out[65]
port 379 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1400 90 0 0 la_data_out[66]
port 380 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1400 90 0 0 la_data_out[67]
port 381 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1400 90 0 0 la_data_out[68]
port 382 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1400 90 0 0 la_data_out[69]
port 383 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1400 90 0 0 la_data_out[6]
port 384 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1400 90 0 0 la_data_out[70]
port 385 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1400 90 0 0 la_data_out[71]
port 386 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1400 90 0 0 la_data_out[72]
port 387 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1400 90 0 0 la_data_out[73]
port 388 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1400 90 0 0 la_data_out[74]
port 389 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1400 90 0 0 la_data_out[75]
port 390 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1400 90 0 0 la_data_out[76]
port 391 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1400 90 0 0 la_data_out[77]
port 392 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1400 90 0 0 la_data_out[78]
port 393 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1400 90 0 0 la_data_out[79]
port 394 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1400 90 0 0 la_data_out[7]
port 395 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1400 90 0 0 la_data_out[80]
port 396 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1400 90 0 0 la_data_out[81]
port 397 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1400 90 0 0 la_data_out[82]
port 398 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1400 90 0 0 la_data_out[83]
port 399 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1400 90 0 0 la_data_out[84]
port 400 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1400 90 0 0 la_data_out[85]
port 401 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1400 90 0 0 la_data_out[86]
port 402 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1400 90 0 0 la_data_out[87]
port 403 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1400 90 0 0 la_data_out[88]
port 404 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1400 90 0 0 la_data_out[89]
port 405 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1400 90 0 0 la_data_out[8]
port 406 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1400 90 0 0 la_data_out[90]
port 407 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1400 90 0 0 la_data_out[91]
port 408 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1400 90 0 0 la_data_out[92]
port 409 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1400 90 0 0 la_data_out[93]
port 410 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1400 90 0 0 la_data_out[94]
port 411 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1400 90 0 0 la_data_out[95]
port 412 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1400 90 0 0 la_data_out[96]
port 413 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1400 90 0 0 la_data_out[97]
port 414 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1400 90 0 0 la_data_out[98]
port 415 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1400 90 0 0 la_data_out[99]
port 416 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1400 90 0 0 la_data_out[9]
port 417 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1400 90 0 0 la_oenb[0]
port 418 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1400 90 0 0 la_oenb[100]
port 419 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1400 90 0 0 la_oenb[101]
port 420 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1400 90 0 0 la_oenb[102]
port 421 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1400 90 0 0 la_oenb[103]
port 422 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1400 90 0 0 la_oenb[104]
port 423 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1400 90 0 0 la_oenb[105]
port 424 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1400 90 0 0 la_oenb[106]
port 425 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1400 90 0 0 la_oenb[107]
port 426 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1400 90 0 0 la_oenb[108]
port 427 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1400 90 0 0 la_oenb[109]
port 428 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1400 90 0 0 la_oenb[10]
port 429 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1400 90 0 0 la_oenb[110]
port 430 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1400 90 0 0 la_oenb[111]
port 431 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1400 90 0 0 la_oenb[112]
port 432 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1400 90 0 0 la_oenb[113]
port 433 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1400 90 0 0 la_oenb[114]
port 434 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1400 90 0 0 la_oenb[115]
port 435 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1400 90 0 0 la_oenb[116]
port 436 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1400 90 0 0 la_oenb[117]
port 437 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1400 90 0 0 la_oenb[118]
port 438 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1400 90 0 0 la_oenb[119]
port 439 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1400 90 0 0 la_oenb[11]
port 440 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1400 90 0 0 la_oenb[120]
port 441 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1400 90 0 0 la_oenb[121]
port 442 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1400 90 0 0 la_oenb[122]
port 443 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1400 90 0 0 la_oenb[123]
port 444 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1400 90 0 0 la_oenb[124]
port 445 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1400 90 0 0 la_oenb[125]
port 446 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1400 90 0 0 la_oenb[126]
port 447 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1400 90 0 0 la_oenb[127]
port 448 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1400 90 0 0 la_oenb[12]
port 449 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1400 90 0 0 la_oenb[13]
port 450 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1400 90 0 0 la_oenb[14]
port 451 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1400 90 0 0 la_oenb[15]
port 452 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1400 90 0 0 la_oenb[16]
port 453 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1400 90 0 0 la_oenb[17]
port 454 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1400 90 0 0 la_oenb[18]
port 455 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1400 90 0 0 la_oenb[19]
port 456 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1400 90 0 0 la_oenb[1]
port 457 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1400 90 0 0 la_oenb[20]
port 458 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1400 90 0 0 la_oenb[21]
port 459 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1400 90 0 0 la_oenb[22]
port 460 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1400 90 0 0 la_oenb[23]
port 461 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1400 90 0 0 la_oenb[24]
port 462 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1400 90 0 0 la_oenb[25]
port 463 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1400 90 0 0 la_oenb[26]
port 464 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1400 90 0 0 la_oenb[27]
port 465 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1400 90 0 0 la_oenb[28]
port 466 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1400 90 0 0 la_oenb[29]
port 467 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1400 90 0 0 la_oenb[2]
port 468 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1400 90 0 0 la_oenb[30]
port 469 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1400 90 0 0 la_oenb[31]
port 470 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1400 90 0 0 la_oenb[32]
port 471 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1400 90 0 0 la_oenb[33]
port 472 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1400 90 0 0 la_oenb[34]
port 473 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1400 90 0 0 la_oenb[35]
port 474 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1400 90 0 0 la_oenb[36]
port 475 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1400 90 0 0 la_oenb[37]
port 476 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1400 90 0 0 la_oenb[38]
port 477 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1400 90 0 0 la_oenb[39]
port 478 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1400 90 0 0 la_oenb[3]
port 479 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1400 90 0 0 la_oenb[40]
port 480 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1400 90 0 0 la_oenb[41]
port 481 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1400 90 0 0 la_oenb[42]
port 482 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1400 90 0 0 la_oenb[43]
port 483 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1400 90 0 0 la_oenb[44]
port 484 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1400 90 0 0 la_oenb[45]
port 485 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1400 90 0 0 la_oenb[46]
port 486 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1400 90 0 0 la_oenb[47]
port 487 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1400 90 0 0 la_oenb[48]
port 488 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1400 90 0 0 la_oenb[49]
port 489 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1400 90 0 0 la_oenb[4]
port 490 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1400 90 0 0 la_oenb[50]
port 491 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1400 90 0 0 la_oenb[51]
port 492 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1400 90 0 0 la_oenb[52]
port 493 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1400 90 0 0 la_oenb[53]
port 494 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1400 90 0 0 la_oenb[54]
port 495 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1400 90 0 0 la_oenb[55]
port 496 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1400 90 0 0 la_oenb[56]
port 497 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1400 90 0 0 la_oenb[57]
port 498 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1400 90 0 0 la_oenb[58]
port 499 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1400 90 0 0 la_oenb[59]
port 500 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1400 90 0 0 la_oenb[5]
port 501 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1400 90 0 0 la_oenb[60]
port 502 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1400 90 0 0 la_oenb[61]
port 503 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1400 90 0 0 la_oenb[62]
port 504 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1400 90 0 0 la_oenb[63]
port 505 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1400 90 0 0 la_oenb[64]
port 506 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1400 90 0 0 la_oenb[65]
port 507 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1400 90 0 0 la_oenb[66]
port 508 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1400 90 0 0 la_oenb[67]
port 509 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1400 90 0 0 la_oenb[68]
port 510 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1400 90 0 0 la_oenb[69]
port 511 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1400 90 0 0 la_oenb[6]
port 512 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1400 90 0 0 la_oenb[70]
port 513 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1400 90 0 0 la_oenb[71]
port 514 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1400 90 0 0 la_oenb[72]
port 515 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1400 90 0 0 la_oenb[73]
port 516 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1400 90 0 0 la_oenb[74]
port 517 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1400 90 0 0 la_oenb[75]
port 518 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1400 90 0 0 la_oenb[76]
port 519 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1400 90 0 0 la_oenb[77]
port 520 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1400 90 0 0 la_oenb[78]
port 521 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1400 90 0 0 la_oenb[79]
port 522 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1400 90 0 0 la_oenb[7]
port 523 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1400 90 0 0 la_oenb[80]
port 524 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1400 90 0 0 la_oenb[81]
port 525 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1400 90 0 0 la_oenb[82]
port 526 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1400 90 0 0 la_oenb[83]
port 527 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1400 90 0 0 la_oenb[84]
port 528 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1400 90 0 0 la_oenb[85]
port 529 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1400 90 0 0 la_oenb[86]
port 530 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1400 90 0 0 la_oenb[87]
port 531 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1400 90 0 0 la_oenb[88]
port 532 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1400 90 0 0 la_oenb[89]
port 533 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1400 90 0 0 la_oenb[8]
port 534 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1400 90 0 0 la_oenb[90]
port 535 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1400 90 0 0 la_oenb[91]
port 536 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1400 90 0 0 la_oenb[92]
port 537 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1400 90 0 0 la_oenb[93]
port 538 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1400 90 0 0 la_oenb[94]
port 539 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1400 90 0 0 la_oenb[95]
port 540 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1400 90 0 0 la_oenb[96]
port 541 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1400 90 0 0 la_oenb[97]
port 542 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1400 90 0 0 la_oenb[98]
port 543 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1400 90 0 0 la_oenb[99]
port 544 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1400 90 0 0 la_oenb[9]
port 545 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1400 90 0 0 user_clock2
port 546 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1400 90 0 0 user_irq[0]
port 547 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1400 90 0 0 user_irq[1]
port 548 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1400 90 0 0 user_irq[2]
port 549 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 1400 90 0 0 wb_clk_i
port 558 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1400 90 0 0 wb_rst_i
port 559 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1400 90 0 0 wbs_ack_o
port 560 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1400 90 0 0 wbs_adr_i[0]
port 561 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1400 90 0 0 wbs_adr_i[10]
port 562 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1400 90 0 0 wbs_adr_i[11]
port 563 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1400 90 0 0 wbs_adr_i[12]
port 564 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1400 90 0 0 wbs_adr_i[13]
port 565 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1400 90 0 0 wbs_adr_i[14]
port 566 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1400 90 0 0 wbs_adr_i[15]
port 567 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1400 90 0 0 wbs_adr_i[16]
port 568 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1400 90 0 0 wbs_adr_i[17]
port 569 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1400 90 0 0 wbs_adr_i[18]
port 570 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1400 90 0 0 wbs_adr_i[19]
port 571 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1400 90 0 0 wbs_adr_i[1]
port 572 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1400 90 0 0 wbs_adr_i[20]
port 573 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1400 90 0 0 wbs_adr_i[21]
port 574 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1400 90 0 0 wbs_adr_i[22]
port 575 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1400 90 0 0 wbs_adr_i[23]
port 576 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1400 90 0 0 wbs_adr_i[24]
port 577 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1400 90 0 0 wbs_adr_i[25]
port 578 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1400 90 0 0 wbs_adr_i[26]
port 579 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1400 90 0 0 wbs_adr_i[27]
port 580 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1400 90 0 0 wbs_adr_i[28]
port 581 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1400 90 0 0 wbs_adr_i[29]
port 582 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1400 90 0 0 wbs_adr_i[2]
port 583 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1400 90 0 0 wbs_adr_i[30]
port 584 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1400 90 0 0 wbs_adr_i[31]
port 585 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1400 90 0 0 wbs_adr_i[3]
port 586 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1400 90 0 0 wbs_adr_i[4]
port 587 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1400 90 0 0 wbs_adr_i[5]
port 588 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1400 90 0 0 wbs_adr_i[6]
port 589 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1400 90 0 0 wbs_adr_i[7]
port 590 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1400 90 0 0 wbs_adr_i[8]
port 591 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1400 90 0 0 wbs_adr_i[9]
port 592 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1400 90 0 0 wbs_cyc_i
port 593 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1400 90 0 0 wbs_dat_i[0]
port 594 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1400 90 0 0 wbs_dat_i[10]
port 595 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1400 90 0 0 wbs_dat_i[11]
port 596 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1400 90 0 0 wbs_dat_i[12]
port 597 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1400 90 0 0 wbs_dat_i[13]
port 598 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1400 90 0 0 wbs_dat_i[14]
port 599 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1400 90 0 0 wbs_dat_i[15]
port 600 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1400 90 0 0 wbs_dat_i[16]
port 601 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1400 90 0 0 wbs_dat_i[17]
port 602 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1400 90 0 0 wbs_dat_i[18]
port 603 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1400 90 0 0 wbs_dat_i[19]
port 604 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1400 90 0 0 wbs_dat_i[1]
port 605 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1400 90 0 0 wbs_dat_i[20]
port 606 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1400 90 0 0 wbs_dat_i[21]
port 607 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1400 90 0 0 wbs_dat_i[22]
port 608 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1400 90 0 0 wbs_dat_i[23]
port 609 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1400 90 0 0 wbs_dat_i[24]
port 610 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1400 90 0 0 wbs_dat_i[25]
port 611 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1400 90 0 0 wbs_dat_i[26]
port 612 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1400 90 0 0 wbs_dat_i[27]
port 613 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1400 90 0 0 wbs_dat_i[28]
port 614 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1400 90 0 0 wbs_dat_i[29]
port 615 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1400 90 0 0 wbs_dat_i[2]
port 616 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1400 90 0 0 wbs_dat_i[30]
port 617 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1400 90 0 0 wbs_dat_i[31]
port 618 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1400 90 0 0 wbs_dat_i[3]
port 619 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1400 90 0 0 wbs_dat_i[4]
port 620 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1400 90 0 0 wbs_dat_i[5]
port 621 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1400 90 0 0 wbs_dat_i[6]
port 622 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1400 90 0 0 wbs_dat_i[7]
port 623 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1400 90 0 0 wbs_dat_i[8]
port 624 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1400 90 0 0 wbs_dat_i[9]
port 625 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1400 90 0 0 wbs_dat_o[0]
port 626 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1400 90 0 0 wbs_dat_o[10]
port 627 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1400 90 0 0 wbs_dat_o[11]
port 628 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1400 90 0 0 wbs_dat_o[12]
port 629 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1400 90 0 0 wbs_dat_o[13]
port 630 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1400 90 0 0 wbs_dat_o[14]
port 631 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1400 90 0 0 wbs_dat_o[15]
port 632 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1400 90 0 0 wbs_dat_o[16]
port 633 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1400 90 0 0 wbs_dat_o[17]
port 634 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1400 90 0 0 wbs_dat_o[18]
port 635 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1400 90 0 0 wbs_dat_o[19]
port 636 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1400 90 0 0 wbs_dat_o[1]
port 637 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1400 90 0 0 wbs_dat_o[20]
port 638 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1400 90 0 0 wbs_dat_o[21]
port 639 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1400 90 0 0 wbs_dat_o[22]
port 640 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1400 90 0 0 wbs_dat_o[23]
port 641 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1400 90 0 0 wbs_dat_o[24]
port 642 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1400 90 0 0 wbs_dat_o[25]
port 643 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1400 90 0 0 wbs_dat_o[26]
port 644 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1400 90 0 0 wbs_dat_o[27]
port 645 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1400 90 0 0 wbs_dat_o[28]
port 646 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1400 90 0 0 wbs_dat_o[29]
port 647 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1400 90 0 0 wbs_dat_o[2]
port 648 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1400 90 0 0 wbs_dat_o[30]
port 649 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1400 90 0 0 wbs_dat_o[31]
port 650 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1400 90 0 0 wbs_dat_o[3]
port 651 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1400 90 0 0 wbs_dat_o[4]
port 652 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1400 90 0 0 wbs_dat_o[5]
port 653 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1400 90 0 0 wbs_dat_o[6]
port 654 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1400 90 0 0 wbs_dat_o[7]
port 655 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1400 90 0 0 wbs_dat_o[8]
port 656 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1400 90 0 0 wbs_dat_o[9]
port 657 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1400 90 0 0 wbs_sel_i[0]
port 658 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1400 90 0 0 wbs_sel_i[1]
port 659 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1400 90 0 0 wbs_sel_i[2]
port 660 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1400 90 0 0 wbs_sel_i[3]
port 661 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1400 90 0 0 wbs_stb_i
port 662 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1400 90 0 0 wbs_we_i
port 663 nsew
flabel metal1 148648 55790 148848 55990 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFET_3V_1nf_1/GSense_nFET_3VD_3Vg_1nf_0.VD_H
flabel metal1 150348 55790 150548 55990 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFET_3V_1nf_1/GSense_nFET_3VD_3Vg_1nf_0.VLow_Src
flabel metal1 149548 55090 149748 55290 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFET_3V_1nf_1/GSense_nFET_3VD_3Vg_1nf_0.VG_H
flabel metal1 60098 145780 60298 145980 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_pfet_1p8Vd_1p8Vg_0/GSense_pFET_1p8VD_1p8Vg_1nf_0.VLow_Src
flabel metal1 58698 145780 58898 145980 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_pfet_1p8Vd_1p8Vg_0/GSense_pFET_1p8VD_1p8Vg_1nf_0.VD_H
flabel metal1 59298 145180 59498 145380 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_pfet_1p8Vd_1p8Vg_0/GSense_pFET_1p8VD_1p8Vg_1nf_0.VG_H
flabel metal1 59238 56578 59438 56778 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_2.GSense_nFET_1f1WL150n_V1_0/VG_H
flabel metal1 60358 55780 60558 55980 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_2.GSense_nFET_1f1WL150n_V1_0.VLow_Src
flabel metal1 58158 55780 58358 55980 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_2.GSense_nFET_1f1WL150n_V1_0.VD_H
flabel metal1 59238 55000 59438 55200 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_2.GSense_nFET_1f1WL150n_V1_0.VG_H
flabel metal1 148658 145340 148858 145540 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_pFET_10Vd_5p5Vg_1nf_0/GSense_pFET_10VD_5Vg_1nf_0.VD_H
flabel metal1 150258 145340 150458 145540 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_pFET_10Vd_5p5Vg_1nf_0/GSense_pFET_10VD_5Vg_1nf_0.VLow_Src
flabel metal1 149458 144640 149658 144840 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_pFET_10Vd_5p5Vg_1nf_0/GSense_pFET_10VD_5Vg_1nf_0.VG_H
flabel metal1 238658 55500 238858 55700 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFT_g5_10Vd_1nf_0/GSense_nFET_10VD_5Vg_1nf_0.VD_H
flabel metal1 239558 54700 239758 54900 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFT_g5_10Vd_1nf_0/GSense_nFET_10VD_5Vg_1nf_0.VG_H
flabel metal1 240358 55500 240558 55700 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFT_g5_10Vd_1nf_0/GSense_nFET_10VD_5Vg_1nf_0.VLow_Src
flabel metal1 239238 146578 239438 146778 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_0.GSense_nFET_1f1WL150n_V1_0/VG_H
flabel metal1 240358 145780 240558 145980 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_0.GSense_nFET_1f1WL150n_V1_0.VLow_Src
flabel metal1 238158 145780 238358 145980 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_0.GSense_nFET_1f1WL150n_V1_0.VD_H
flabel metal1 239238 145000 239438 145200 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_0.GSense_nFET_1f1WL150n_V1_0.VG_H
flabel metal1 330098 145780 330298 145980 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_pfet_1p8Vd_1p8Vg_1/GSense_pFET_1p8VD_1p8Vg_1nf_0.VLow_Src
flabel metal1 328698 145780 328898 145980 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_pfet_1p8Vd_1p8Vg_1/GSense_pFET_1p8VD_1p8Vg_1nf_0.VD_H
flabel metal1 329298 145180 329498 145380 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_pfet_1p8Vd_1p8Vg_1/GSense_pFET_1p8VD_1p8Vg_1nf_0.VG_H
flabel metal1 329238 56578 329438 56778 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_1.GSense_nFET_1f1WL150n_V1_0/VG_H
flabel metal1 330358 55780 330558 55980 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_1.GSense_nFET_1f1WL150n_V1_0.VLow_Src
flabel metal1 328158 55780 328358 55980 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_1.GSense_nFET_1f1WL150n_V1_0.VD_H
flabel metal1 329238 55000 329438 55200 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_1.GSense_nFET_1f1WL150n_V1_0.VG_H
flabel metal1 418648 55790 418848 55990 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFET_3V_1nf_0/GSense_nFET_3VD_3Vg_1nf_0.VD_H
flabel metal1 420348 55790 420548 55990 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFET_3V_1nf_0/GSense_nFET_3VD_3Vg_1nf_0.VLow_Src
flabel metal1 419548 55090 419748 55290 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFET_3V_1nf_0/GSense_nFET_3VD_3Vg_1nf_0.VG_H
flabel metal1 418658 145340 418858 145540 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_pFET_10Vd_5p5Vg_1nf_1/GSense_pFET_10VD_5Vg_1nf_0.VD_H
flabel metal1 420258 145340 420458 145540 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_pFET_10Vd_5p5Vg_1nf_1/GSense_pFET_10VD_5Vg_1nf_0.VLow_Src
flabel metal1 419458 144640 419658 144840 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_pFET_10Vd_5p5Vg_1nf_1/GSense_pFET_10VD_5Vg_1nf_0.VG_H
flabel metal1 508658 55500 508858 55700 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFT_g5_10Vd_1nf_1/GSense_nFET_10VD_5Vg_1nf_0.VD_H
flabel metal1 509558 54700 509758 54900 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFT_g5_10Vd_1nf_1/GSense_nFET_10VD_5Vg_1nf_0.VG_H
flabel metal1 510358 55500 510558 55700 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFT_g5_10Vd_1nf_1/GSense_nFET_10VD_5Vg_1nf_0.VLow_Src
flabel metal1 509238 146578 509438 146778 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_3.GSense_nFET_1f1WL150n_V1_0/VG_H
flabel metal1 510358 145780 510558 145980 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_3.GSense_nFET_1f1WL150n_V1_0.VLow_Src
flabel metal1 508158 145780 508358 145980 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_3.GSense_nFET_1f1WL150n_V1_0.VD_H
flabel metal1 509238 145000 509438 145200 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_3.GSense_nFET_1f1WL150n_V1_0.VG_H
flabel metal1 58723 251816 58923 252016 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_3p3V_5nF_Contacts_V2_0/GSense_nFET_3VD_3Vg_5nf_V2_1.VD_H
flabel metal1 58873 250866 59073 251066 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_3p3V_5nF_Contacts_V2_0/GSense_nFET_3VD_3Vg_5nf_V2_1.VG_H
flabel metal1 60073 251816 60273 252016 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_3p3V_5nF_Contacts_V2_0/GSense_nFET_3VD_3Vg_5nf_V2_1.VLow_Src
flabel metal1 148628 250704 148828 250904 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_10nF_Contacts_0/GSense_nFET_3VD_3Vg_10nf_V2_0.VG_H
flabel metal1 147088 251430 147288 251630 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_10nF_Contacts_0/GSense_nFET_3VD_3Vg_10nf_V2_0.VD_H
flabel metal1 151792 251414 151992 251614 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_10nF_Contacts_0/GSense_nFET_3VD_3Vg_10nf_V2_0.VLow_Src
flabel metal1 238210 250500 238410 250700 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3p3Vd_3VG_51NF_LTherm_Contacts_0/GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH_0.VG_H
flabel metal1 232726 251690 232926 251890 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3p3Vd_3VG_51NF_LTherm_Contacts_0/GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH_0.VD_H
flabel metal1 249570 251616 249770 251816 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3p3Vd_3VG_51NF_LTherm_Contacts_0/GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH_0.VLow_Src
flabel metal1 326649 249619 326849 249819 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50nF_Therm_FET12_0/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Mid_Therm_0.VG_H
flabel metal1 321165 250809 321365 251009 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50nF_Therm_FET12_0/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Mid_Therm_0.VD_H
flabel metal1 338009 250735 338209 250935 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50nF_Therm_FET12_0/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Mid_Therm_0.VLow_Src
flabel metal1 417292 250215 417492 250415 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_0/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0.VG_H
flabel metal1 411808 251405 412008 251605 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_0/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0.VD_H
flabel metal1 428652 251331 428852 251531 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_0/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0.VLow_Src
flabel metal1 507292 250215 507492 250415 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_1/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0.VG_H
flabel metal1 501808 251405 502008 251605 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_1/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0.VD_H
flabel metal1 518652 251331 518852 251531 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_1/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0.VLow_Src
flabel metal1 57292 370215 57492 370415 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_2/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0.VG_H
flabel metal1 51808 371405 52008 371605 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_2/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0.VD_H
flabel metal1 68652 371331 68852 371531 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_2/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0.VLow_Src
flabel metal1 147292 370215 147492 370415 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_5/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0.VG_H
flabel metal1 141808 371405 142008 371605 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_5/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0.VD_H
flabel metal1 158652 371331 158852 371531 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_5/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0.VLow_Src
flabel metal1 236649 369619 236849 369819 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50nF_Therm_FET12_3/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Mid_Therm_0.VG_H
flabel metal1 231165 370809 231365 371009 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50nF_Therm_FET12_3/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Mid_Therm_0.VD_H
flabel metal1 248009 370735 248209 370935 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50nF_Therm_FET12_3/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Mid_Therm_0.VLow_Src
flabel metal1 327832 370892 328032 371092 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3p3Vd_3VG_51NF_LTherm_Contacts_2/GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH_0.VG_H
flabel metal1 322348 372082 322548 372282 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3p3Vd_3VG_51NF_LTherm_Contacts_2/GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH_0.VD_H
flabel metal1 339192 372008 339392 372208 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3p3Vd_3VG_51NF_LTherm_Contacts_2/GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH_0.VLow_Src
flabel metal1 419504 370908 419704 371108 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_10nF_Contacts_2/GSense_nFET_3VD_3Vg_10nf_V2_0.VG_H
flabel metal1 417964 371634 418164 371834 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_10nF_Contacts_2/GSense_nFET_3VD_3Vg_10nf_V2_0.VD_H
flabel metal1 422668 371618 422868 371818 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_10nF_Contacts_2/GSense_nFET_3VD_3Vg_10nf_V2_0.VLow_Src
flabel metal1 508723 371816 508923 372016 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_3p3V_5nF_Contacts_V2_1/GSense_nFET_3VD_3Vg_5nf_V2_1.VD_H
flabel metal1 508873 370866 509073 371066 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_3p3V_5nF_Contacts_V2_1/GSense_nFET_3VD_3Vg_5nf_V2_1.VG_H
flabel metal1 510073 371816 510273 372016 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_3p3V_5nF_Contacts_V2_1/GSense_nFET_3VD_3Vg_5nf_V2_1.VLow_Src
flabel metal1 59504 490908 59704 491108 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_10nF_Contacts_3/GSense_nFET_3VD_3Vg_10nf_V2_0.VG_H
flabel metal1 57964 491634 58164 491834 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_10nF_Contacts_3/GSense_nFET_3VD_3Vg_10nf_V2_0.VD_H
flabel metal1 62668 491618 62868 491818 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_10nF_Contacts_3/GSense_nFET_3VD_3Vg_10nf_V2_0.VLow_Src
flabel metal1 147292 490215 147492 490415 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_3/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0.VG_H
flabel metal1 141808 491405 142008 491605 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_3/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0.VD_H
flabel metal1 158652 491331 158852 491531 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_3/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0.VLow_Src
flabel metal1 236649 489619 236849 489819 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50nF_Therm_FET12_1/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Mid_Therm_0.VG_H
flabel metal1 231165 490809 231365 491009 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50nF_Therm_FET12_1/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Mid_Therm_0.VD_H
flabel metal1 248009 490735 248209 490935 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_50nF_Therm_FET12_1/GSense_nFET_3VD_3Vg_51nf_V2AllGates_Mid_Therm_0.VLow_Src
flabel metal1 327832 490892 328032 491092 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3p3Vd_3VG_51NF_LTherm_Contacts_1/GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH_0.VG_H
flabel metal1 322348 492082 322548 492282 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3p3Vd_3VG_51NF_LTherm_Contacts_1/GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH_0.VD_H
flabel metal1 339192 492008 339392 492208 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3p3Vd_3VG_51NF_LTherm_Contacts_1/GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH_0.VLow_Src
flabel metal1 418723 491816 418923 492016 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_3p3V_5nF_Contacts_V2_2/GSense_nFET_3VD_3Vg_5nf_V2_1.VD_H
flabel metal1 418873 490866 419073 491066 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_3p3V_5nF_Contacts_V2_2/GSense_nFET_3VD_3Vg_5nf_V2_1.VG_H
flabel metal1 420073 491816 420273 492016 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_3p3V_5nF_Contacts_V2_2/GSense_nFET_3VD_3Vg_5nf_V2_1.VLow_Src
flabel metal1 509504 490908 509704 491108 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_10nF_Contacts_1/GSense_nFET_3VD_3Vg_10nf_V2_0.VG_H
flabel metal1 507964 491634 508164 491834 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_10nF_Contacts_1/GSense_nFET_3VD_3Vg_10nf_V2_0.VD_H
flabel metal1 512668 491618 512868 491818 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/nFET_3VD_3VG_10nF_Contacts_1/GSense_nFET_3VD_3Vg_10nf_V2_0.VLow_Src
flabel metal1 58648 580790 58848 580990 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFET_3V_1nf_2/GSense_nFET_3VD_3Vg_1nf_0.VD_H
flabel metal1 60348 580790 60548 580990 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFET_3V_1nf_2/GSense_nFET_3VD_3Vg_1nf_0.VLow_Src
flabel metal1 59548 580090 59748 580290 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFET_3V_1nf_2/GSense_nFET_3VD_3Vg_1nf_0.VG_H
flabel metal1 148658 580500 148858 580700 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFT_g5_10Vd_1nf_2/GSense_nFET_10VD_5Vg_1nf_0.VD_H
flabel metal1 149558 579700 149758 579900 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFT_g5_10Vd_1nf_2/GSense_nFET_10VD_5Vg_1nf_0.VG_H
flabel metal1 150358 580500 150558 580700 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFT_g5_10Vd_1nf_2/GSense_nFET_10VD_5Vg_1nf_0.VLow_Src
flabel metal1 239238 581578 239438 581778 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_4.GSense_nFET_1f1WL150n_V1_0/VG_H
flabel metal1 240358 580780 240558 580980 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_4.GSense_nFET_1f1WL150n_V1_0.VLow_Src
flabel metal1 238158 580780 238358 580980 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_4.GSense_nFET_1f1WL150n_V1_0.VD_H
flabel metal1 239238 580000 239438 580200 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_4.GSense_nFET_1f1WL150n_V1_0.VG_H
flabel metal1 328658 580340 328858 580540 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_pFET_10Vd_5p5Vg_1nf_2/GSense_pFET_10VD_5Vg_1nf_0.VD_H
flabel metal1 330258 580340 330458 580540 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_pFET_10Vd_5p5Vg_1nf_2/GSense_pFET_10VD_5Vg_1nf_0.VLow_Src
flabel metal1 329458 579640 329658 579840 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_pFET_10Vd_5p5Vg_1nf_2/GSense_pFET_10VD_5Vg_1nf_0.VG_H
flabel metal1 58648 655790 58848 655990 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFET_3V_1nf_3/GSense_nFET_3VD_3Vg_1nf_0.VD_H
flabel metal1 60348 655790 60548 655990 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFET_3V_1nf_3/GSense_nFET_3VD_3Vg_1nf_0.VLow_Src
flabel metal1 59548 655090 59748 655290 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_nFET_3V_1nf_3/GSense_nFET_3VD_3Vg_1nf_0.VG_H
flabel metal1 149238 656578 149438 656778 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_5.GSense_nFET_1f1WL150n_V1_0/VG_H
flabel metal1 150358 655780 150558 655980 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_5.GSense_nFET_1f1WL150n_V1_0.VLow_Src
flabel metal1 148158 655780 148358 655980 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_5.GSense_nFET_1f1WL150n_V1_0.VD_H
flabel metal1 149238 655000 149438 655200 0 FreeSans 256 0 0 0 transistor_layout_20240603_0/GSense_nFET_1W015L_1F_Contacts_5.GSense_nFET_1f1WL150n_V1_0.VG_H
flabel metal1 240098 655780 240298 655980 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_pfet_1p8Vd_1p8Vg_2/GSense_pFET_1p8VD_1p8Vg_1nf_0.VLow_Src
flabel metal1 238698 655780 238898 655980 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_pfet_1p8Vd_1p8Vg_2/GSense_pFET_1p8VD_1p8Vg_1nf_0.VD_H
flabel metal1 239298 655180 239498 655380 0 FreeSans 160 0 0 0 transistor_layout_20240603_0/GSense_Contacts_pfet_1p8Vd_1p8Vg_2/GSense_pFET_1p8VD_1p8Vg_1nf_0.VG_H
flabel metal1 418460 657264 418660 657464 0 FreeSans 160 0 0 0 GSense_pFET_10Vd_5p5Vg_1nf_1/GSense_pFET_10VD_5Vg_1nf_0.VD_H
flabel metal1 420060 657264 420260 657464 0 FreeSans 160 0 0 0 GSense_pFET_10Vd_5p5Vg_1nf_1/GSense_pFET_10VD_5Vg_1nf_0.VLow_Src
flabel metal1 419260 656564 419460 656764 0 FreeSans 160 0 0 0 GSense_pFET_10Vd_5p5Vg_1nf_1/GSense_pFET_10VD_5Vg_1nf_0.VG_H
flabel metal1 509040 658502 509240 658702 0 FreeSans 256 0 0 0 GSense_nFET_1W015L_1F_Contacts_3.GSense_nFET_1f1WL150n_V1_0/VG_H
flabel metal1 510160 657704 510360 657904 0 FreeSans 256 0 0 0 GSense_nFET_1W015L_1F_Contacts_3.GSense_nFET_1f1WL150n_V1_0.VLow_Src
flabel metal1 507960 657704 508160 657904 0 FreeSans 256 0 0 0 GSense_nFET_1W015L_1F_Contacts_3.GSense_nFET_1f1WL150n_V1_0.VD_H
flabel metal1 509040 656924 509240 657124 0 FreeSans 256 0 0 0 GSense_nFET_1W015L_1F_Contacts_3.GSense_nFET_1f1WL150n_V1_0.VG_H
flabel metal1 329040 658502 329240 658702 0 FreeSans 256 0 0 0 GSense_nFET_1W015L_1F_Contacts_1.GSense_nFET_1f1WL150n_V1_0/VG_H
flabel metal1 330160 657704 330360 657904 0 FreeSans 256 0 0 0 GSense_nFET_1W015L_1F_Contacts_1.GSense_nFET_1f1WL150n_V1_0.VLow_Src
flabel metal1 327960 657704 328160 657904 0 FreeSans 256 0 0 0 GSense_nFET_1W015L_1F_Contacts_1.GSense_nFET_1f1WL150n_V1_0.VD_H
flabel metal1 329040 656924 329240 657124 0 FreeSans 256 0 0 0 GSense_nFET_1W015L_1F_Contacts_1.GSense_nFET_1f1WL150n_V1_0.VG_H
flabel metal1 508460 582424 508660 582624 0 FreeSans 256 0 0 0 GSense_Contacts_nFT_g5_10Vd_1nf_1/GSense_nFET_10VD_5Vg_1nf_0.VD_H
flabel metal1 509360 581624 509560 581824 0 FreeSans 256 0 0 0 GSense_Contacts_nFT_g5_10Vd_1nf_1/GSense_nFET_10VD_5Vg_1nf_0.VG_H
flabel metal1 510160 582424 510360 582624 0 FreeSans 256 0 0 0 GSense_Contacts_nFT_g5_10Vd_1nf_1/GSense_nFET_10VD_5Vg_1nf_0.VLow_Src
flabel metal1 418450 582714 418650 582914 0 FreeSans 160 0 0 0 GSense_Contacts_nFET_3V_1nf_0/GSense_nFET_3VD_3Vg_1nf_0.VD_H
flabel metal1 420150 582714 420350 582914 0 FreeSans 160 0 0 0 GSense_Contacts_nFET_3V_1nf_0/GSense_nFET_3VD_3Vg_1nf_0.VLow_Src
flabel metal1 419350 582014 419550 582214 0 FreeSans 160 0 0 0 GSense_Contacts_nFET_3V_1nf_0/GSense_nFET_3VD_3Vg_1nf_0.VG_H
<< end >>
