magic
tech sky130A
magscale 1 2
timestamp 1717253661
<< metal1 >>
rect 2690 -222 2830 -204
rect 2768 -336 2830 -222
rect 2690 -356 2830 -336
<< via1 >>
rect 2690 -336 2768 -222
<< metal2 >>
rect 852 4928 1112 4968
rect 852 4712 900 4928
rect 1062 4712 1112 4928
rect 852 2368 1112 4712
rect 2814 -204 3259 -202
rect 2690 -222 3259 -204
rect 2768 -336 3259 -222
rect 2690 -356 3259 -336
rect 3413 -356 3430 -202
rect -880 -2622 -712 -2232
rect -880 -2774 -852 -2622
rect -738 -2774 -712 -2622
rect -880 -2802 -712 -2774
<< via2 >>
rect 900 4712 1062 4928
rect 3259 -356 3413 -202
rect -852 -2774 -738 -2622
<< metal3 >>
rect 512 8122 1420 8264
rect 512 7716 738 8122
rect 1220 7716 1420 8122
rect 512 6024 1420 7716
rect 838 4928 1088 6024
rect 838 4712 900 4928
rect 1062 4712 1088 4928
rect 838 4664 1088 4712
rect -2564 -840 -1332 -82
rect 3254 -202 3418 -197
rect 3254 -356 3259 -202
rect 3413 -319 4577 -202
rect 5373 -319 6247 -299
rect 3413 -356 6247 -319
rect 3254 -361 3418 -356
rect 4423 -600 6247 -356
rect -2564 -1040 -2514 -840
rect -2314 -1040 -1090 -840
rect 4423 -885 5550 -600
rect -2564 -1390 -1332 -1040
rect 4419 -1050 5550 -885
rect 6000 -1050 6247 -600
rect 4419 -1335 6247 -1050
rect -882 -2622 -710 -2570
rect -882 -2774 -852 -2622
rect -738 -2774 -710 -2622
rect 430 -2640 662 -2232
rect 430 -2680 672 -2640
rect -882 -2996 -710 -2774
rect -1268 -5270 -386 -2996
rect 420 -2998 672 -2680
rect -1268 -5884 -1046 -5270
rect -522 -5884 -386 -5270
rect -1268 -6080 -386 -5884
rect 24 -5252 962 -2998
rect 24 -5900 274 -5252
rect 788 -5900 962 -5252
rect 24 -6094 962 -5900
<< via3 >>
rect 738 7716 1220 8122
rect -2514 -1040 -2314 -840
rect 5550 -1050 6000 -600
rect -1046 -5884 -522 -5270
rect 274 -5900 788 -5252
<< metal4 >>
rect 520 13418 1470 13660
rect 520 12936 722 13418
rect 1300 12936 1470 13418
rect 520 8122 1470 12936
rect 520 7716 738 8122
rect 1220 7716 1470 8122
rect 520 7476 1470 7716
rect -5238 -780 -2276 -82
rect -5238 -1100 -5204 -780
rect -4884 -840 -2276 -780
rect -4884 -1040 -2514 -840
rect -2314 -1040 -2276 -840
rect -4884 -1100 -2276 -1040
rect -5238 -1408 -2276 -1100
rect 5344 -185 8884 -100
rect 5344 -316 8893 -185
rect 5344 -600 8168 -316
rect 5344 -1050 5550 -600
rect 6000 -950 8168 -600
rect 8820 -950 8893 -316
rect 6000 -1050 8893 -950
rect 5344 -1061 8893 -1050
rect 5344 -1370 8884 -1061
rect -1276 -5270 -384 -4546
rect 24 -5242 980 -4556
rect 2402 -5242 3352 -5214
rect -1276 -5884 -1046 -5270
rect -522 -5884 -384 -5270
rect -1276 -7950 -384 -5884
rect 8 -5252 3352 -5242
rect 8 -5900 274 -5252
rect 788 -5900 3352 -5252
rect 8 -6116 3352 -5900
rect -1276 -9076 -1166 -7950
rect -522 -9076 -384 -7950
rect -1276 -9188 -384 -9076
rect 2402 -7928 3352 -6116
rect 2402 -9072 2586 -7928
rect 3188 -9072 3352 -7928
rect 2402 -9548 3352 -9072
<< via4 >>
rect 722 12936 1300 13418
rect -5204 -1100 -4884 -780
rect 8168 -950 8820 -316
rect -1166 -9076 -522 -7950
rect 2586 -9072 3188 -7928
<< metal5 >>
rect -28066 17000 -12066 25780
rect -28200 16982 0 17000
rect -28200 16000 1512 16982
rect -28066 9580 -12066 16000
rect -762 15998 1512 16000
rect 394 13418 1512 15998
rect 394 12936 722 13418
rect 1300 12936 1512 13418
rect 394 12666 1512 12936
rect -28000 -86 -12000 7100
rect 15030 54 31030 7066
rect -28000 -90 -4910 -86
rect -28000 -780 -4852 -90
rect -28000 -1100 -5204 -780
rect -4884 -1100 -4852 -780
rect -28000 -1376 -4852 -1100
rect 8000 -316 31030 54
rect 8000 -950 8168 -316
rect 8820 -950 31030 -316
rect -28000 -9100 -12000 -1376
rect 8000 -1486 31030 -950
rect -1334 -7950 -366 -7354
rect -1334 -9076 -1166 -7950
rect -522 -9076 -366 -7950
rect -28080 -19776 -12080 -11622
rect -1334 -19776 -366 -9076
rect 2366 -7928 3376 -7352
rect 2366 -9072 2586 -7928
rect 3188 -9072 3376 -7928
rect 2366 -19612 3376 -9072
rect 15030 -9134 31030 -1486
rect 2332 -19628 5378 -19612
rect 15030 -19628 31030 -11764
rect -28080 -20702 -326 -19776
rect -28080 -27822 -12080 -20702
rect 2332 -20744 31030 -19628
rect 15002 -20852 31030 -20744
rect 15030 -27964 31030 -20852
<< glass >>
rect -27600 9800 -12466 25380
rect -27600 -8700 -12400 6700
rect 15430 -8734 30630 6666
rect -27680 -27400 -12480 -12020
rect 15430 -27564 30630 -12164
<< end >>
