magic
tech sky130A
timestamp 1717370063
<< pwell >>
rect -2114 -150 2114 150
<< nnmos >>
rect -2000 -21 -1950 21
rect -1921 -21 -1871 21
rect -1842 -21 -1792 21
rect -1763 -21 -1713 21
rect -1684 -21 -1634 21
rect -1605 -21 -1555 21
rect -1526 -21 -1476 21
rect -1447 -21 -1397 21
rect -1368 -21 -1318 21
rect -1289 -21 -1239 21
rect -1210 -21 -1160 21
rect -1131 -21 -1081 21
rect -1052 -21 -1002 21
rect -973 -21 -923 21
rect -894 -21 -844 21
rect -815 -21 -765 21
rect -736 -21 -686 21
rect -657 -21 -607 21
rect -578 -21 -528 21
rect -499 -21 -449 21
rect -420 -21 -370 21
rect -341 -21 -291 21
rect -262 -21 -212 21
rect -183 -21 -133 21
rect -104 -21 -54 21
rect -25 -21 25 21
rect 54 -21 104 21
rect 133 -21 183 21
rect 212 -21 262 21
rect 291 -21 341 21
rect 370 -21 420 21
rect 449 -21 499 21
rect 528 -21 578 21
rect 607 -21 657 21
rect 686 -21 736 21
rect 765 -21 815 21
rect 844 -21 894 21
rect 923 -21 973 21
rect 1002 -21 1052 21
rect 1081 -21 1131 21
rect 1160 -21 1210 21
rect 1239 -21 1289 21
rect 1318 -21 1368 21
rect 1397 -21 1447 21
rect 1476 -21 1526 21
rect 1555 -21 1605 21
rect 1634 -21 1684 21
rect 1713 -21 1763 21
rect 1792 -21 1842 21
rect 1871 -21 1921 21
rect 1950 -21 2000 21
<< mvndiff >>
rect -2029 15 -2000 21
rect -2029 -15 -2023 15
rect -2006 -15 -2000 15
rect -2029 -21 -2000 -15
rect -1950 15 -1921 21
rect -1950 -15 -1944 15
rect -1927 -15 -1921 15
rect -1950 -21 -1921 -15
rect -1871 15 -1842 21
rect -1871 -15 -1865 15
rect -1848 -15 -1842 15
rect -1871 -21 -1842 -15
rect -1792 15 -1763 21
rect -1792 -15 -1786 15
rect -1769 -15 -1763 15
rect -1792 -21 -1763 -15
rect -1713 15 -1684 21
rect -1713 -15 -1707 15
rect -1690 -15 -1684 15
rect -1713 -21 -1684 -15
rect -1634 15 -1605 21
rect -1634 -15 -1628 15
rect -1611 -15 -1605 15
rect -1634 -21 -1605 -15
rect -1555 15 -1526 21
rect -1555 -15 -1549 15
rect -1532 -15 -1526 15
rect -1555 -21 -1526 -15
rect -1476 15 -1447 21
rect -1476 -15 -1470 15
rect -1453 -15 -1447 15
rect -1476 -21 -1447 -15
rect -1397 15 -1368 21
rect -1397 -15 -1391 15
rect -1374 -15 -1368 15
rect -1397 -21 -1368 -15
rect -1318 15 -1289 21
rect -1318 -15 -1312 15
rect -1295 -15 -1289 15
rect -1318 -21 -1289 -15
rect -1239 15 -1210 21
rect -1239 -15 -1233 15
rect -1216 -15 -1210 15
rect -1239 -21 -1210 -15
rect -1160 15 -1131 21
rect -1160 -15 -1154 15
rect -1137 -15 -1131 15
rect -1160 -21 -1131 -15
rect -1081 15 -1052 21
rect -1081 -15 -1075 15
rect -1058 -15 -1052 15
rect -1081 -21 -1052 -15
rect -1002 15 -973 21
rect -1002 -15 -996 15
rect -979 -15 -973 15
rect -1002 -21 -973 -15
rect -923 15 -894 21
rect -923 -15 -917 15
rect -900 -15 -894 15
rect -923 -21 -894 -15
rect -844 15 -815 21
rect -844 -15 -838 15
rect -821 -15 -815 15
rect -844 -21 -815 -15
rect -765 15 -736 21
rect -765 -15 -759 15
rect -742 -15 -736 15
rect -765 -21 -736 -15
rect -686 15 -657 21
rect -686 -15 -680 15
rect -663 -15 -657 15
rect -686 -21 -657 -15
rect -607 15 -578 21
rect -607 -15 -601 15
rect -584 -15 -578 15
rect -607 -21 -578 -15
rect -528 15 -499 21
rect -528 -15 -522 15
rect -505 -15 -499 15
rect -528 -21 -499 -15
rect -449 15 -420 21
rect -449 -15 -443 15
rect -426 -15 -420 15
rect -449 -21 -420 -15
rect -370 15 -341 21
rect -370 -15 -364 15
rect -347 -15 -341 15
rect -370 -21 -341 -15
rect -291 15 -262 21
rect -291 -15 -285 15
rect -268 -15 -262 15
rect -291 -21 -262 -15
rect -212 15 -183 21
rect -212 -15 -206 15
rect -189 -15 -183 15
rect -212 -21 -183 -15
rect -133 15 -104 21
rect -133 -15 -127 15
rect -110 -15 -104 15
rect -133 -21 -104 -15
rect -54 15 -25 21
rect -54 -15 -48 15
rect -31 -15 -25 15
rect -54 -21 -25 -15
rect 25 15 54 21
rect 25 -15 31 15
rect 48 -15 54 15
rect 25 -21 54 -15
rect 104 15 133 21
rect 104 -15 110 15
rect 127 -15 133 15
rect 104 -21 133 -15
rect 183 15 212 21
rect 183 -15 189 15
rect 206 -15 212 15
rect 183 -21 212 -15
rect 262 15 291 21
rect 262 -15 268 15
rect 285 -15 291 15
rect 262 -21 291 -15
rect 341 15 370 21
rect 341 -15 347 15
rect 364 -15 370 15
rect 341 -21 370 -15
rect 420 15 449 21
rect 420 -15 426 15
rect 443 -15 449 15
rect 420 -21 449 -15
rect 499 15 528 21
rect 499 -15 505 15
rect 522 -15 528 15
rect 499 -21 528 -15
rect 578 15 607 21
rect 578 -15 584 15
rect 601 -15 607 15
rect 578 -21 607 -15
rect 657 15 686 21
rect 657 -15 663 15
rect 680 -15 686 15
rect 657 -21 686 -15
rect 736 15 765 21
rect 736 -15 742 15
rect 759 -15 765 15
rect 736 -21 765 -15
rect 815 15 844 21
rect 815 -15 821 15
rect 838 -15 844 15
rect 815 -21 844 -15
rect 894 15 923 21
rect 894 -15 900 15
rect 917 -15 923 15
rect 894 -21 923 -15
rect 973 15 1002 21
rect 973 -15 979 15
rect 996 -15 1002 15
rect 973 -21 1002 -15
rect 1052 15 1081 21
rect 1052 -15 1058 15
rect 1075 -15 1081 15
rect 1052 -21 1081 -15
rect 1131 15 1160 21
rect 1131 -15 1137 15
rect 1154 -15 1160 15
rect 1131 -21 1160 -15
rect 1210 15 1239 21
rect 1210 -15 1216 15
rect 1233 -15 1239 15
rect 1210 -21 1239 -15
rect 1289 15 1318 21
rect 1289 -15 1295 15
rect 1312 -15 1318 15
rect 1289 -21 1318 -15
rect 1368 15 1397 21
rect 1368 -15 1374 15
rect 1391 -15 1397 15
rect 1368 -21 1397 -15
rect 1447 15 1476 21
rect 1447 -15 1453 15
rect 1470 -15 1476 15
rect 1447 -21 1476 -15
rect 1526 15 1555 21
rect 1526 -15 1532 15
rect 1549 -15 1555 15
rect 1526 -21 1555 -15
rect 1605 15 1634 21
rect 1605 -15 1611 15
rect 1628 -15 1634 15
rect 1605 -21 1634 -15
rect 1684 15 1713 21
rect 1684 -15 1690 15
rect 1707 -15 1713 15
rect 1684 -21 1713 -15
rect 1763 15 1792 21
rect 1763 -15 1769 15
rect 1786 -15 1792 15
rect 1763 -21 1792 -15
rect 1842 15 1871 21
rect 1842 -15 1848 15
rect 1865 -15 1871 15
rect 1842 -21 1871 -15
rect 1921 15 1950 21
rect 1921 -15 1927 15
rect 1944 -15 1950 15
rect 1921 -21 1950 -15
rect 2000 15 2029 21
rect 2000 -15 2006 15
rect 2023 -15 2029 15
rect 2000 -21 2029 -15
<< mvndiffc >>
rect -2023 -15 -2006 15
rect -1944 -15 -1927 15
rect -1865 -15 -1848 15
rect -1786 -15 -1769 15
rect -1707 -15 -1690 15
rect -1628 -15 -1611 15
rect -1549 -15 -1532 15
rect -1470 -15 -1453 15
rect -1391 -15 -1374 15
rect -1312 -15 -1295 15
rect -1233 -15 -1216 15
rect -1154 -15 -1137 15
rect -1075 -15 -1058 15
rect -996 -15 -979 15
rect -917 -15 -900 15
rect -838 -15 -821 15
rect -759 -15 -742 15
rect -680 -15 -663 15
rect -601 -15 -584 15
rect -522 -15 -505 15
rect -443 -15 -426 15
rect -364 -15 -347 15
rect -285 -15 -268 15
rect -206 -15 -189 15
rect -127 -15 -110 15
rect -48 -15 -31 15
rect 31 -15 48 15
rect 110 -15 127 15
rect 189 -15 206 15
rect 268 -15 285 15
rect 347 -15 364 15
rect 426 -15 443 15
rect 505 -15 522 15
rect 584 -15 601 15
rect 663 -15 680 15
rect 742 -15 759 15
rect 821 -15 838 15
rect 900 -15 917 15
rect 979 -15 996 15
rect 1058 -15 1075 15
rect 1137 -15 1154 15
rect 1216 -15 1233 15
rect 1295 -15 1312 15
rect 1374 -15 1391 15
rect 1453 -15 1470 15
rect 1532 -15 1549 15
rect 1611 -15 1628 15
rect 1690 -15 1707 15
rect 1769 -15 1786 15
rect 1848 -15 1865 15
rect 1927 -15 1944 15
rect 2006 -15 2023 15
<< mvpsubdiff >>
rect -2096 126 2096 132
rect -2096 109 -2042 126
rect 2042 109 2096 126
rect -2096 103 2096 109
rect -2096 78 -2067 103
rect -2096 -78 -2090 78
rect -2073 -78 -2067 78
rect 2067 78 2096 103
rect -2096 -103 -2067 -78
rect 2067 -78 2073 78
rect 2090 -78 2096 78
rect 2067 -103 2096 -78
rect -2096 -109 2096 -103
rect -2096 -126 -2042 -109
rect 2042 -126 2096 -109
rect -2096 -132 2096 -126
<< mvpsubdiffcont >>
rect -2042 109 2042 126
rect -2090 -78 -2073 78
rect 2073 -78 2090 78
rect -2042 -126 2042 -109
<< poly >>
rect -2000 57 -1950 65
rect -2000 40 -1992 57
rect -1958 40 -1950 57
rect -2000 21 -1950 40
rect -1921 57 -1871 65
rect -1921 40 -1913 57
rect -1879 40 -1871 57
rect -1921 21 -1871 40
rect -1842 57 -1792 65
rect -1842 40 -1834 57
rect -1800 40 -1792 57
rect -1842 21 -1792 40
rect -1763 57 -1713 65
rect -1763 40 -1755 57
rect -1721 40 -1713 57
rect -1763 21 -1713 40
rect -1684 57 -1634 65
rect -1684 40 -1676 57
rect -1642 40 -1634 57
rect -1684 21 -1634 40
rect -1605 57 -1555 65
rect -1605 40 -1597 57
rect -1563 40 -1555 57
rect -1605 21 -1555 40
rect -1526 57 -1476 65
rect -1526 40 -1518 57
rect -1484 40 -1476 57
rect -1526 21 -1476 40
rect -1447 57 -1397 65
rect -1447 40 -1439 57
rect -1405 40 -1397 57
rect -1447 21 -1397 40
rect -1368 57 -1318 65
rect -1368 40 -1360 57
rect -1326 40 -1318 57
rect -1368 21 -1318 40
rect -1289 57 -1239 65
rect -1289 40 -1281 57
rect -1247 40 -1239 57
rect -1289 21 -1239 40
rect -1210 57 -1160 65
rect -1210 40 -1202 57
rect -1168 40 -1160 57
rect -1210 21 -1160 40
rect -1131 57 -1081 65
rect -1131 40 -1123 57
rect -1089 40 -1081 57
rect -1131 21 -1081 40
rect -1052 57 -1002 65
rect -1052 40 -1044 57
rect -1010 40 -1002 57
rect -1052 21 -1002 40
rect -973 57 -923 65
rect -973 40 -965 57
rect -931 40 -923 57
rect -973 21 -923 40
rect -894 57 -844 65
rect -894 40 -886 57
rect -852 40 -844 57
rect -894 21 -844 40
rect -815 57 -765 65
rect -815 40 -807 57
rect -773 40 -765 57
rect -815 21 -765 40
rect -736 57 -686 65
rect -736 40 -728 57
rect -694 40 -686 57
rect -736 21 -686 40
rect -657 57 -607 65
rect -657 40 -649 57
rect -615 40 -607 57
rect -657 21 -607 40
rect -578 57 -528 65
rect -578 40 -570 57
rect -536 40 -528 57
rect -578 21 -528 40
rect -499 57 -449 65
rect -499 40 -491 57
rect -457 40 -449 57
rect -499 21 -449 40
rect -420 57 -370 65
rect -420 40 -412 57
rect -378 40 -370 57
rect -420 21 -370 40
rect -341 57 -291 65
rect -341 40 -333 57
rect -299 40 -291 57
rect -341 21 -291 40
rect -262 57 -212 65
rect -262 40 -254 57
rect -220 40 -212 57
rect -262 21 -212 40
rect -183 57 -133 65
rect -183 40 -175 57
rect -141 40 -133 57
rect -183 21 -133 40
rect -104 57 -54 65
rect -104 40 -96 57
rect -62 40 -54 57
rect -104 21 -54 40
rect -25 57 25 65
rect -25 40 -17 57
rect 17 40 25 57
rect -25 21 25 40
rect 54 57 104 65
rect 54 40 62 57
rect 96 40 104 57
rect 54 21 104 40
rect 133 57 183 65
rect 133 40 141 57
rect 175 40 183 57
rect 133 21 183 40
rect 212 57 262 65
rect 212 40 220 57
rect 254 40 262 57
rect 212 21 262 40
rect 291 57 341 65
rect 291 40 299 57
rect 333 40 341 57
rect 291 21 341 40
rect 370 57 420 65
rect 370 40 378 57
rect 412 40 420 57
rect 370 21 420 40
rect 449 57 499 65
rect 449 40 457 57
rect 491 40 499 57
rect 449 21 499 40
rect 528 57 578 65
rect 528 40 536 57
rect 570 40 578 57
rect 528 21 578 40
rect 607 57 657 65
rect 607 40 615 57
rect 649 40 657 57
rect 607 21 657 40
rect 686 57 736 65
rect 686 40 694 57
rect 728 40 736 57
rect 686 21 736 40
rect 765 57 815 65
rect 765 40 773 57
rect 807 40 815 57
rect 765 21 815 40
rect 844 57 894 65
rect 844 40 852 57
rect 886 40 894 57
rect 844 21 894 40
rect 923 57 973 65
rect 923 40 931 57
rect 965 40 973 57
rect 923 21 973 40
rect 1002 57 1052 65
rect 1002 40 1010 57
rect 1044 40 1052 57
rect 1002 21 1052 40
rect 1081 57 1131 65
rect 1081 40 1089 57
rect 1123 40 1131 57
rect 1081 21 1131 40
rect 1160 57 1210 65
rect 1160 40 1168 57
rect 1202 40 1210 57
rect 1160 21 1210 40
rect 1239 57 1289 65
rect 1239 40 1247 57
rect 1281 40 1289 57
rect 1239 21 1289 40
rect 1318 57 1368 65
rect 1318 40 1326 57
rect 1360 40 1368 57
rect 1318 21 1368 40
rect 1397 57 1447 65
rect 1397 40 1405 57
rect 1439 40 1447 57
rect 1397 21 1447 40
rect 1476 57 1526 65
rect 1476 40 1484 57
rect 1518 40 1526 57
rect 1476 21 1526 40
rect 1555 57 1605 65
rect 1555 40 1563 57
rect 1597 40 1605 57
rect 1555 21 1605 40
rect 1634 57 1684 65
rect 1634 40 1642 57
rect 1676 40 1684 57
rect 1634 21 1684 40
rect 1713 57 1763 65
rect 1713 40 1721 57
rect 1755 40 1763 57
rect 1713 21 1763 40
rect 1792 57 1842 65
rect 1792 40 1800 57
rect 1834 40 1842 57
rect 1792 21 1842 40
rect 1871 57 1921 65
rect 1871 40 1879 57
rect 1913 40 1921 57
rect 1871 21 1921 40
rect 1950 57 2000 65
rect 1950 40 1958 57
rect 1992 40 2000 57
rect 1950 21 2000 40
rect -2000 -40 -1950 -21
rect -2000 -57 -1992 -40
rect -1958 -57 -1950 -40
rect -2000 -65 -1950 -57
rect -1921 -40 -1871 -21
rect -1921 -57 -1913 -40
rect -1879 -57 -1871 -40
rect -1921 -65 -1871 -57
rect -1842 -40 -1792 -21
rect -1842 -57 -1834 -40
rect -1800 -57 -1792 -40
rect -1842 -65 -1792 -57
rect -1763 -40 -1713 -21
rect -1763 -57 -1755 -40
rect -1721 -57 -1713 -40
rect -1763 -65 -1713 -57
rect -1684 -40 -1634 -21
rect -1684 -57 -1676 -40
rect -1642 -57 -1634 -40
rect -1684 -65 -1634 -57
rect -1605 -40 -1555 -21
rect -1605 -57 -1597 -40
rect -1563 -57 -1555 -40
rect -1605 -65 -1555 -57
rect -1526 -40 -1476 -21
rect -1526 -57 -1518 -40
rect -1484 -57 -1476 -40
rect -1526 -65 -1476 -57
rect -1447 -40 -1397 -21
rect -1447 -57 -1439 -40
rect -1405 -57 -1397 -40
rect -1447 -65 -1397 -57
rect -1368 -40 -1318 -21
rect -1368 -57 -1360 -40
rect -1326 -57 -1318 -40
rect -1368 -65 -1318 -57
rect -1289 -40 -1239 -21
rect -1289 -57 -1281 -40
rect -1247 -57 -1239 -40
rect -1289 -65 -1239 -57
rect -1210 -40 -1160 -21
rect -1210 -57 -1202 -40
rect -1168 -57 -1160 -40
rect -1210 -65 -1160 -57
rect -1131 -40 -1081 -21
rect -1131 -57 -1123 -40
rect -1089 -57 -1081 -40
rect -1131 -65 -1081 -57
rect -1052 -40 -1002 -21
rect -1052 -57 -1044 -40
rect -1010 -57 -1002 -40
rect -1052 -65 -1002 -57
rect -973 -40 -923 -21
rect -973 -57 -965 -40
rect -931 -57 -923 -40
rect -973 -65 -923 -57
rect -894 -40 -844 -21
rect -894 -57 -886 -40
rect -852 -57 -844 -40
rect -894 -65 -844 -57
rect -815 -40 -765 -21
rect -815 -57 -807 -40
rect -773 -57 -765 -40
rect -815 -65 -765 -57
rect -736 -40 -686 -21
rect -736 -57 -728 -40
rect -694 -57 -686 -40
rect -736 -65 -686 -57
rect -657 -40 -607 -21
rect -657 -57 -649 -40
rect -615 -57 -607 -40
rect -657 -65 -607 -57
rect -578 -40 -528 -21
rect -578 -57 -570 -40
rect -536 -57 -528 -40
rect -578 -65 -528 -57
rect -499 -40 -449 -21
rect -499 -57 -491 -40
rect -457 -57 -449 -40
rect -499 -65 -449 -57
rect -420 -40 -370 -21
rect -420 -57 -412 -40
rect -378 -57 -370 -40
rect -420 -65 -370 -57
rect -341 -40 -291 -21
rect -341 -57 -333 -40
rect -299 -57 -291 -40
rect -341 -65 -291 -57
rect -262 -40 -212 -21
rect -262 -57 -254 -40
rect -220 -57 -212 -40
rect -262 -65 -212 -57
rect -183 -40 -133 -21
rect -183 -57 -175 -40
rect -141 -57 -133 -40
rect -183 -65 -133 -57
rect -104 -40 -54 -21
rect -104 -57 -96 -40
rect -62 -57 -54 -40
rect -104 -65 -54 -57
rect -25 -40 25 -21
rect -25 -57 -17 -40
rect 17 -57 25 -40
rect -25 -65 25 -57
rect 54 -40 104 -21
rect 54 -57 62 -40
rect 96 -57 104 -40
rect 54 -65 104 -57
rect 133 -40 183 -21
rect 133 -57 141 -40
rect 175 -57 183 -40
rect 133 -65 183 -57
rect 212 -40 262 -21
rect 212 -57 220 -40
rect 254 -57 262 -40
rect 212 -65 262 -57
rect 291 -40 341 -21
rect 291 -57 299 -40
rect 333 -57 341 -40
rect 291 -65 341 -57
rect 370 -40 420 -21
rect 370 -57 378 -40
rect 412 -57 420 -40
rect 370 -65 420 -57
rect 449 -40 499 -21
rect 449 -57 457 -40
rect 491 -57 499 -40
rect 449 -65 499 -57
rect 528 -40 578 -21
rect 528 -57 536 -40
rect 570 -57 578 -40
rect 528 -65 578 -57
rect 607 -40 657 -21
rect 607 -57 615 -40
rect 649 -57 657 -40
rect 607 -65 657 -57
rect 686 -40 736 -21
rect 686 -57 694 -40
rect 728 -57 736 -40
rect 686 -65 736 -57
rect 765 -40 815 -21
rect 765 -57 773 -40
rect 807 -57 815 -40
rect 765 -65 815 -57
rect 844 -40 894 -21
rect 844 -57 852 -40
rect 886 -57 894 -40
rect 844 -65 894 -57
rect 923 -40 973 -21
rect 923 -57 931 -40
rect 965 -57 973 -40
rect 923 -65 973 -57
rect 1002 -40 1052 -21
rect 1002 -57 1010 -40
rect 1044 -57 1052 -40
rect 1002 -65 1052 -57
rect 1081 -40 1131 -21
rect 1081 -57 1089 -40
rect 1123 -57 1131 -40
rect 1081 -65 1131 -57
rect 1160 -40 1210 -21
rect 1160 -57 1168 -40
rect 1202 -57 1210 -40
rect 1160 -65 1210 -57
rect 1239 -40 1289 -21
rect 1239 -57 1247 -40
rect 1281 -57 1289 -40
rect 1239 -65 1289 -57
rect 1318 -40 1368 -21
rect 1318 -57 1326 -40
rect 1360 -57 1368 -40
rect 1318 -65 1368 -57
rect 1397 -40 1447 -21
rect 1397 -57 1405 -40
rect 1439 -57 1447 -40
rect 1397 -65 1447 -57
rect 1476 -40 1526 -21
rect 1476 -57 1484 -40
rect 1518 -57 1526 -40
rect 1476 -65 1526 -57
rect 1555 -40 1605 -21
rect 1555 -57 1563 -40
rect 1597 -57 1605 -40
rect 1555 -65 1605 -57
rect 1634 -40 1684 -21
rect 1634 -57 1642 -40
rect 1676 -57 1684 -40
rect 1634 -65 1684 -57
rect 1713 -40 1763 -21
rect 1713 -57 1721 -40
rect 1755 -57 1763 -40
rect 1713 -65 1763 -57
rect 1792 -40 1842 -21
rect 1792 -57 1800 -40
rect 1834 -57 1842 -40
rect 1792 -65 1842 -57
rect 1871 -40 1921 -21
rect 1871 -57 1879 -40
rect 1913 -57 1921 -40
rect 1871 -65 1921 -57
rect 1950 -40 2000 -21
rect 1950 -57 1958 -40
rect 1992 -57 2000 -40
rect 1950 -65 2000 -57
<< polycont >>
rect -1992 40 -1958 57
rect -1913 40 -1879 57
rect -1834 40 -1800 57
rect -1755 40 -1721 57
rect -1676 40 -1642 57
rect -1597 40 -1563 57
rect -1518 40 -1484 57
rect -1439 40 -1405 57
rect -1360 40 -1326 57
rect -1281 40 -1247 57
rect -1202 40 -1168 57
rect -1123 40 -1089 57
rect -1044 40 -1010 57
rect -965 40 -931 57
rect -886 40 -852 57
rect -807 40 -773 57
rect -728 40 -694 57
rect -649 40 -615 57
rect -570 40 -536 57
rect -491 40 -457 57
rect -412 40 -378 57
rect -333 40 -299 57
rect -254 40 -220 57
rect -175 40 -141 57
rect -96 40 -62 57
rect -17 40 17 57
rect 62 40 96 57
rect 141 40 175 57
rect 220 40 254 57
rect 299 40 333 57
rect 378 40 412 57
rect 457 40 491 57
rect 536 40 570 57
rect 615 40 649 57
rect 694 40 728 57
rect 773 40 807 57
rect 852 40 886 57
rect 931 40 965 57
rect 1010 40 1044 57
rect 1089 40 1123 57
rect 1168 40 1202 57
rect 1247 40 1281 57
rect 1326 40 1360 57
rect 1405 40 1439 57
rect 1484 40 1518 57
rect 1563 40 1597 57
rect 1642 40 1676 57
rect 1721 40 1755 57
rect 1800 40 1834 57
rect 1879 40 1913 57
rect 1958 40 1992 57
rect -1992 -57 -1958 -40
rect -1913 -57 -1879 -40
rect -1834 -57 -1800 -40
rect -1755 -57 -1721 -40
rect -1676 -57 -1642 -40
rect -1597 -57 -1563 -40
rect -1518 -57 -1484 -40
rect -1439 -57 -1405 -40
rect -1360 -57 -1326 -40
rect -1281 -57 -1247 -40
rect -1202 -57 -1168 -40
rect -1123 -57 -1089 -40
rect -1044 -57 -1010 -40
rect -965 -57 -931 -40
rect -886 -57 -852 -40
rect -807 -57 -773 -40
rect -728 -57 -694 -40
rect -649 -57 -615 -40
rect -570 -57 -536 -40
rect -491 -57 -457 -40
rect -412 -57 -378 -40
rect -333 -57 -299 -40
rect -254 -57 -220 -40
rect -175 -57 -141 -40
rect -96 -57 -62 -40
rect -17 -57 17 -40
rect 62 -57 96 -40
rect 141 -57 175 -40
rect 220 -57 254 -40
rect 299 -57 333 -40
rect 378 -57 412 -40
rect 457 -57 491 -40
rect 536 -57 570 -40
rect 615 -57 649 -40
rect 694 -57 728 -40
rect 773 -57 807 -40
rect 852 -57 886 -40
rect 931 -57 965 -40
rect 1010 -57 1044 -40
rect 1089 -57 1123 -40
rect 1168 -57 1202 -40
rect 1247 -57 1281 -40
rect 1326 -57 1360 -40
rect 1405 -57 1439 -40
rect 1484 -57 1518 -40
rect 1563 -57 1597 -40
rect 1642 -57 1676 -40
rect 1721 -57 1755 -40
rect 1800 -57 1834 -40
rect 1879 -57 1913 -40
rect 1958 -57 1992 -40
<< locali >>
rect -2090 109 -2042 126
rect 2042 109 2090 126
rect -2090 78 -2073 109
rect 2073 78 2090 109
rect -2000 40 -1992 57
rect -1958 40 -1950 57
rect -1921 40 -1913 57
rect -1879 40 -1871 57
rect -1842 40 -1834 57
rect -1800 40 -1792 57
rect -1763 40 -1755 57
rect -1721 40 -1713 57
rect -1684 40 -1676 57
rect -1642 40 -1634 57
rect -1605 40 -1597 57
rect -1563 40 -1555 57
rect -1526 40 -1518 57
rect -1484 40 -1476 57
rect -1447 40 -1439 57
rect -1405 40 -1397 57
rect -1368 40 -1360 57
rect -1326 40 -1318 57
rect -1289 40 -1281 57
rect -1247 40 -1239 57
rect -1210 40 -1202 57
rect -1168 40 -1160 57
rect -1131 40 -1123 57
rect -1089 40 -1081 57
rect -1052 40 -1044 57
rect -1010 40 -1002 57
rect -973 40 -965 57
rect -931 40 -923 57
rect -894 40 -886 57
rect -852 40 -844 57
rect -815 40 -807 57
rect -773 40 -765 57
rect -736 40 -728 57
rect -694 40 -686 57
rect -657 40 -649 57
rect -615 40 -607 57
rect -578 40 -570 57
rect -536 40 -528 57
rect -499 40 -491 57
rect -457 40 -449 57
rect -420 40 -412 57
rect -378 40 -370 57
rect -341 40 -333 57
rect -299 40 -291 57
rect -262 40 -254 57
rect -220 40 -212 57
rect -183 40 -175 57
rect -141 40 -133 57
rect -104 40 -96 57
rect -62 40 -54 57
rect -25 40 -17 57
rect 17 40 25 57
rect 54 40 62 57
rect 96 40 104 57
rect 133 40 141 57
rect 175 40 183 57
rect 212 40 220 57
rect 254 40 262 57
rect 291 40 299 57
rect 333 40 341 57
rect 370 40 378 57
rect 412 40 420 57
rect 449 40 457 57
rect 491 40 499 57
rect 528 40 536 57
rect 570 40 578 57
rect 607 40 615 57
rect 649 40 657 57
rect 686 40 694 57
rect 728 40 736 57
rect 765 40 773 57
rect 807 40 815 57
rect 844 40 852 57
rect 886 40 894 57
rect 923 40 931 57
rect 965 40 973 57
rect 1002 40 1010 57
rect 1044 40 1052 57
rect 1081 40 1089 57
rect 1123 40 1131 57
rect 1160 40 1168 57
rect 1202 40 1210 57
rect 1239 40 1247 57
rect 1281 40 1289 57
rect 1318 40 1326 57
rect 1360 40 1368 57
rect 1397 40 1405 57
rect 1439 40 1447 57
rect 1476 40 1484 57
rect 1518 40 1526 57
rect 1555 40 1563 57
rect 1597 40 1605 57
rect 1634 40 1642 57
rect 1676 40 1684 57
rect 1713 40 1721 57
rect 1755 40 1763 57
rect 1792 40 1800 57
rect 1834 40 1842 57
rect 1871 40 1879 57
rect 1913 40 1921 57
rect 1950 40 1958 57
rect 1992 40 2000 57
rect -2023 15 -2006 23
rect -2023 -23 -2006 -15
rect -1944 15 -1927 23
rect -1944 -23 -1927 -15
rect -1865 15 -1848 23
rect -1865 -23 -1848 -15
rect -1786 15 -1769 23
rect -1786 -23 -1769 -15
rect -1707 15 -1690 23
rect -1707 -23 -1690 -15
rect -1628 15 -1611 23
rect -1628 -23 -1611 -15
rect -1549 15 -1532 23
rect -1549 -23 -1532 -15
rect -1470 15 -1453 23
rect -1470 -23 -1453 -15
rect -1391 15 -1374 23
rect -1391 -23 -1374 -15
rect -1312 15 -1295 23
rect -1312 -23 -1295 -15
rect -1233 15 -1216 23
rect -1233 -23 -1216 -15
rect -1154 15 -1137 23
rect -1154 -23 -1137 -15
rect -1075 15 -1058 23
rect -1075 -23 -1058 -15
rect -996 15 -979 23
rect -996 -23 -979 -15
rect -917 15 -900 23
rect -917 -23 -900 -15
rect -838 15 -821 23
rect -838 -23 -821 -15
rect -759 15 -742 23
rect -759 -23 -742 -15
rect -680 15 -663 23
rect -680 -23 -663 -15
rect -601 15 -584 23
rect -601 -23 -584 -15
rect -522 15 -505 23
rect -522 -23 -505 -15
rect -443 15 -426 23
rect -443 -23 -426 -15
rect -364 15 -347 23
rect -364 -23 -347 -15
rect -285 15 -268 23
rect -285 -23 -268 -15
rect -206 15 -189 23
rect -206 -23 -189 -15
rect -127 15 -110 23
rect -127 -23 -110 -15
rect -48 15 -31 23
rect -48 -23 -31 -15
rect 31 15 48 23
rect 31 -23 48 -15
rect 110 15 127 23
rect 110 -23 127 -15
rect 189 15 206 23
rect 189 -23 206 -15
rect 268 15 285 23
rect 268 -23 285 -15
rect 347 15 364 23
rect 347 -23 364 -15
rect 426 15 443 23
rect 426 -23 443 -15
rect 505 15 522 23
rect 505 -23 522 -15
rect 584 15 601 23
rect 584 -23 601 -15
rect 663 15 680 23
rect 663 -23 680 -15
rect 742 15 759 23
rect 742 -23 759 -15
rect 821 15 838 23
rect 821 -23 838 -15
rect 900 15 917 23
rect 900 -23 917 -15
rect 979 15 996 23
rect 979 -23 996 -15
rect 1058 15 1075 23
rect 1058 -23 1075 -15
rect 1137 15 1154 23
rect 1137 -23 1154 -15
rect 1216 15 1233 23
rect 1216 -23 1233 -15
rect 1295 15 1312 23
rect 1295 -23 1312 -15
rect 1374 15 1391 23
rect 1374 -23 1391 -15
rect 1453 15 1470 23
rect 1453 -23 1470 -15
rect 1532 15 1549 23
rect 1532 -23 1549 -15
rect 1611 15 1628 23
rect 1611 -23 1628 -15
rect 1690 15 1707 23
rect 1690 -23 1707 -15
rect 1769 15 1786 23
rect 1769 -23 1786 -15
rect 1848 15 1865 23
rect 1848 -23 1865 -15
rect 1927 15 1944 23
rect 1927 -23 1944 -15
rect 2006 15 2023 23
rect 2006 -23 2023 -15
rect -2000 -57 -1992 -40
rect -1958 -57 -1950 -40
rect -1921 -57 -1913 -40
rect -1879 -57 -1871 -40
rect -1842 -57 -1834 -40
rect -1800 -57 -1792 -40
rect -1763 -57 -1755 -40
rect -1721 -57 -1713 -40
rect -1684 -57 -1676 -40
rect -1642 -57 -1634 -40
rect -1605 -57 -1597 -40
rect -1563 -57 -1555 -40
rect -1526 -57 -1518 -40
rect -1484 -57 -1476 -40
rect -1447 -57 -1439 -40
rect -1405 -57 -1397 -40
rect -1368 -57 -1360 -40
rect -1326 -57 -1318 -40
rect -1289 -57 -1281 -40
rect -1247 -57 -1239 -40
rect -1210 -57 -1202 -40
rect -1168 -57 -1160 -40
rect -1131 -57 -1123 -40
rect -1089 -57 -1081 -40
rect -1052 -57 -1044 -40
rect -1010 -57 -1002 -40
rect -973 -57 -965 -40
rect -931 -57 -923 -40
rect -894 -57 -886 -40
rect -852 -57 -844 -40
rect -815 -57 -807 -40
rect -773 -57 -765 -40
rect -736 -57 -728 -40
rect -694 -57 -686 -40
rect -657 -57 -649 -40
rect -615 -57 -607 -40
rect -578 -57 -570 -40
rect -536 -57 -528 -40
rect -499 -57 -491 -40
rect -457 -57 -449 -40
rect -420 -57 -412 -40
rect -378 -57 -370 -40
rect -341 -57 -333 -40
rect -299 -57 -291 -40
rect -262 -57 -254 -40
rect -220 -57 -212 -40
rect -183 -57 -175 -40
rect -141 -57 -133 -40
rect -104 -57 -96 -40
rect -62 -57 -54 -40
rect -25 -57 -17 -40
rect 17 -57 25 -40
rect 54 -57 62 -40
rect 96 -57 104 -40
rect 133 -57 141 -40
rect 175 -57 183 -40
rect 212 -57 220 -40
rect 254 -57 262 -40
rect 291 -57 299 -40
rect 333 -57 341 -40
rect 370 -57 378 -40
rect 412 -57 420 -40
rect 449 -57 457 -40
rect 491 -57 499 -40
rect 528 -57 536 -40
rect 570 -57 578 -40
rect 607 -57 615 -40
rect 649 -57 657 -40
rect 686 -57 694 -40
rect 728 -57 736 -40
rect 765 -57 773 -40
rect 807 -57 815 -40
rect 844 -57 852 -40
rect 886 -57 894 -40
rect 923 -57 931 -40
rect 965 -57 973 -40
rect 1002 -57 1010 -40
rect 1044 -57 1052 -40
rect 1081 -57 1089 -40
rect 1123 -57 1131 -40
rect 1160 -57 1168 -40
rect 1202 -57 1210 -40
rect 1239 -57 1247 -40
rect 1281 -57 1289 -40
rect 1318 -57 1326 -40
rect 1360 -57 1368 -40
rect 1397 -57 1405 -40
rect 1439 -57 1447 -40
rect 1476 -57 1484 -40
rect 1518 -57 1526 -40
rect 1555 -57 1563 -40
rect 1597 -57 1605 -40
rect 1634 -57 1642 -40
rect 1676 -57 1684 -40
rect 1713 -57 1721 -40
rect 1755 -57 1763 -40
rect 1792 -57 1800 -40
rect 1834 -57 1842 -40
rect 1871 -57 1879 -40
rect 1913 -57 1921 -40
rect 1950 -57 1958 -40
rect 1992 -57 2000 -40
rect -2090 -109 -2073 -78
rect 2073 -109 2090 -78
rect -2090 -126 -2042 -109
rect 2042 -126 2090 -109
<< viali >>
rect -1992 40 -1958 57
rect -1913 40 -1879 57
rect -1834 40 -1800 57
rect -1755 40 -1721 57
rect -1676 40 -1642 57
rect -1597 40 -1563 57
rect -1518 40 -1484 57
rect -1439 40 -1405 57
rect -1360 40 -1326 57
rect -1281 40 -1247 57
rect -1202 40 -1168 57
rect -1123 40 -1089 57
rect -1044 40 -1010 57
rect -965 40 -931 57
rect -886 40 -852 57
rect -807 40 -773 57
rect -728 40 -694 57
rect -649 40 -615 57
rect -570 40 -536 57
rect -491 40 -457 57
rect -412 40 -378 57
rect -333 40 -299 57
rect -254 40 -220 57
rect -175 40 -141 57
rect -96 40 -62 57
rect -17 40 17 57
rect 62 40 96 57
rect 141 40 175 57
rect 220 40 254 57
rect 299 40 333 57
rect 378 40 412 57
rect 457 40 491 57
rect 536 40 570 57
rect 615 40 649 57
rect 694 40 728 57
rect 773 40 807 57
rect 852 40 886 57
rect 931 40 965 57
rect 1010 40 1044 57
rect 1089 40 1123 57
rect 1168 40 1202 57
rect 1247 40 1281 57
rect 1326 40 1360 57
rect 1405 40 1439 57
rect 1484 40 1518 57
rect 1563 40 1597 57
rect 1642 40 1676 57
rect 1721 40 1755 57
rect 1800 40 1834 57
rect 1879 40 1913 57
rect 1958 40 1992 57
rect -2023 -15 -2006 15
rect -1944 -15 -1927 15
rect -1865 -15 -1848 15
rect -1786 -15 -1769 15
rect -1707 -15 -1690 15
rect -1628 -15 -1611 15
rect -1549 -15 -1532 15
rect -1470 -15 -1453 15
rect -1391 -15 -1374 15
rect -1312 -15 -1295 15
rect -1233 -15 -1216 15
rect -1154 -15 -1137 15
rect -1075 -15 -1058 15
rect -996 -15 -979 15
rect -917 -15 -900 15
rect -838 -15 -821 15
rect -759 -15 -742 15
rect -680 -15 -663 15
rect -601 -15 -584 15
rect -522 -15 -505 15
rect -443 -15 -426 15
rect -364 -15 -347 15
rect -285 -15 -268 15
rect -206 -15 -189 15
rect -127 -15 -110 15
rect -48 -15 -31 15
rect 31 -15 48 15
rect 110 -15 127 15
rect 189 -15 206 15
rect 268 -15 285 15
rect 347 -15 364 15
rect 426 -15 443 15
rect 505 -15 522 15
rect 584 -15 601 15
rect 663 -15 680 15
rect 742 -15 759 15
rect 821 -15 838 15
rect 900 -15 917 15
rect 979 -15 996 15
rect 1058 -15 1075 15
rect 1137 -15 1154 15
rect 1216 -15 1233 15
rect 1295 -15 1312 15
rect 1374 -15 1391 15
rect 1453 -15 1470 15
rect 1532 -15 1549 15
rect 1611 -15 1628 15
rect 1690 -15 1707 15
rect 1769 -15 1786 15
rect 1848 -15 1865 15
rect 1927 -15 1944 15
rect 2006 -15 2023 15
rect -1992 -57 -1958 -40
rect -1913 -57 -1879 -40
rect -1834 -57 -1800 -40
rect -1755 -57 -1721 -40
rect -1676 -57 -1642 -40
rect -1597 -57 -1563 -40
rect -1518 -57 -1484 -40
rect -1439 -57 -1405 -40
rect -1360 -57 -1326 -40
rect -1281 -57 -1247 -40
rect -1202 -57 -1168 -40
rect -1123 -57 -1089 -40
rect -1044 -57 -1010 -40
rect -965 -57 -931 -40
rect -886 -57 -852 -40
rect -807 -57 -773 -40
rect -728 -57 -694 -40
rect -649 -57 -615 -40
rect -570 -57 -536 -40
rect -491 -57 -457 -40
rect -412 -57 -378 -40
rect -333 -57 -299 -40
rect -254 -57 -220 -40
rect -175 -57 -141 -40
rect -96 -57 -62 -40
rect -17 -57 17 -40
rect 62 -57 96 -40
rect 141 -57 175 -40
rect 220 -57 254 -40
rect 299 -57 333 -40
rect 378 -57 412 -40
rect 457 -57 491 -40
rect 536 -57 570 -40
rect 615 -57 649 -40
rect 694 -57 728 -40
rect 773 -57 807 -40
rect 852 -57 886 -40
rect 931 -57 965 -40
rect 1010 -57 1044 -40
rect 1089 -57 1123 -40
rect 1168 -57 1202 -40
rect 1247 -57 1281 -40
rect 1326 -57 1360 -40
rect 1405 -57 1439 -40
rect 1484 -57 1518 -40
rect 1563 -57 1597 -40
rect 1642 -57 1676 -40
rect 1721 -57 1755 -40
rect 1800 -57 1834 -40
rect 1879 -57 1913 -40
rect 1958 -57 1992 -40
<< metal1 >>
rect -1998 57 -1952 60
rect -1998 40 -1992 57
rect -1958 40 -1952 57
rect -1998 37 -1952 40
rect -1919 57 -1873 60
rect -1919 40 -1913 57
rect -1879 40 -1873 57
rect -1919 37 -1873 40
rect -1840 57 -1794 60
rect -1840 40 -1834 57
rect -1800 40 -1794 57
rect -1840 37 -1794 40
rect -1761 57 -1715 60
rect -1761 40 -1755 57
rect -1721 40 -1715 57
rect -1761 37 -1715 40
rect -1682 57 -1636 60
rect -1682 40 -1676 57
rect -1642 40 -1636 57
rect -1682 37 -1636 40
rect -1603 57 -1557 60
rect -1603 40 -1597 57
rect -1563 40 -1557 57
rect -1603 37 -1557 40
rect -1524 57 -1478 60
rect -1524 40 -1518 57
rect -1484 40 -1478 57
rect -1524 37 -1478 40
rect -1445 57 -1399 60
rect -1445 40 -1439 57
rect -1405 40 -1399 57
rect -1445 37 -1399 40
rect -1366 57 -1320 60
rect -1366 40 -1360 57
rect -1326 40 -1320 57
rect -1366 37 -1320 40
rect -1287 57 -1241 60
rect -1287 40 -1281 57
rect -1247 40 -1241 57
rect -1287 37 -1241 40
rect -1208 57 -1162 60
rect -1208 40 -1202 57
rect -1168 40 -1162 57
rect -1208 37 -1162 40
rect -1129 57 -1083 60
rect -1129 40 -1123 57
rect -1089 40 -1083 57
rect -1129 37 -1083 40
rect -1050 57 -1004 60
rect -1050 40 -1044 57
rect -1010 40 -1004 57
rect -1050 37 -1004 40
rect -971 57 -925 60
rect -971 40 -965 57
rect -931 40 -925 57
rect -971 37 -925 40
rect -892 57 -846 60
rect -892 40 -886 57
rect -852 40 -846 57
rect -892 37 -846 40
rect -813 57 -767 60
rect -813 40 -807 57
rect -773 40 -767 57
rect -813 37 -767 40
rect -734 57 -688 60
rect -734 40 -728 57
rect -694 40 -688 57
rect -734 37 -688 40
rect -655 57 -609 60
rect -655 40 -649 57
rect -615 40 -609 57
rect -655 37 -609 40
rect -576 57 -530 60
rect -576 40 -570 57
rect -536 40 -530 57
rect -576 37 -530 40
rect -497 57 -451 60
rect -497 40 -491 57
rect -457 40 -451 57
rect -497 37 -451 40
rect -418 57 -372 60
rect -418 40 -412 57
rect -378 40 -372 57
rect -418 37 -372 40
rect -339 57 -293 60
rect -339 40 -333 57
rect -299 40 -293 57
rect -339 37 -293 40
rect -260 57 -214 60
rect -260 40 -254 57
rect -220 40 -214 57
rect -260 37 -214 40
rect -181 57 -135 60
rect -181 40 -175 57
rect -141 40 -135 57
rect -181 37 -135 40
rect -102 57 -56 60
rect -102 40 -96 57
rect -62 40 -56 57
rect -102 37 -56 40
rect -23 57 23 60
rect -23 40 -17 57
rect 17 40 23 57
rect -23 37 23 40
rect 56 57 102 60
rect 56 40 62 57
rect 96 40 102 57
rect 56 37 102 40
rect 135 57 181 60
rect 135 40 141 57
rect 175 40 181 57
rect 135 37 181 40
rect 214 57 260 60
rect 214 40 220 57
rect 254 40 260 57
rect 214 37 260 40
rect 293 57 339 60
rect 293 40 299 57
rect 333 40 339 57
rect 293 37 339 40
rect 372 57 418 60
rect 372 40 378 57
rect 412 40 418 57
rect 372 37 418 40
rect 451 57 497 60
rect 451 40 457 57
rect 491 40 497 57
rect 451 37 497 40
rect 530 57 576 60
rect 530 40 536 57
rect 570 40 576 57
rect 530 37 576 40
rect 609 57 655 60
rect 609 40 615 57
rect 649 40 655 57
rect 609 37 655 40
rect 688 57 734 60
rect 688 40 694 57
rect 728 40 734 57
rect 688 37 734 40
rect 767 57 813 60
rect 767 40 773 57
rect 807 40 813 57
rect 767 37 813 40
rect 846 57 892 60
rect 846 40 852 57
rect 886 40 892 57
rect 846 37 892 40
rect 925 57 971 60
rect 925 40 931 57
rect 965 40 971 57
rect 925 37 971 40
rect 1004 57 1050 60
rect 1004 40 1010 57
rect 1044 40 1050 57
rect 1004 37 1050 40
rect 1083 57 1129 60
rect 1083 40 1089 57
rect 1123 40 1129 57
rect 1083 37 1129 40
rect 1162 57 1208 60
rect 1162 40 1168 57
rect 1202 40 1208 57
rect 1162 37 1208 40
rect 1241 57 1287 60
rect 1241 40 1247 57
rect 1281 40 1287 57
rect 1241 37 1287 40
rect 1320 57 1366 60
rect 1320 40 1326 57
rect 1360 40 1366 57
rect 1320 37 1366 40
rect 1399 57 1445 60
rect 1399 40 1405 57
rect 1439 40 1445 57
rect 1399 37 1445 40
rect 1478 57 1524 60
rect 1478 40 1484 57
rect 1518 40 1524 57
rect 1478 37 1524 40
rect 1557 57 1603 60
rect 1557 40 1563 57
rect 1597 40 1603 57
rect 1557 37 1603 40
rect 1636 57 1682 60
rect 1636 40 1642 57
rect 1676 40 1682 57
rect 1636 37 1682 40
rect 1715 57 1761 60
rect 1715 40 1721 57
rect 1755 40 1761 57
rect 1715 37 1761 40
rect 1794 57 1840 60
rect 1794 40 1800 57
rect 1834 40 1840 57
rect 1794 37 1840 40
rect 1873 57 1919 60
rect 1873 40 1879 57
rect 1913 40 1919 57
rect 1873 37 1919 40
rect 1952 57 1998 60
rect 1952 40 1958 57
rect 1992 40 1998 57
rect 1952 37 1998 40
rect -2026 15 -2003 21
rect -2026 -15 -2023 15
rect -2006 -15 -2003 15
rect -2026 -21 -2003 -15
rect -1947 15 -1924 21
rect -1947 -15 -1944 15
rect -1927 -15 -1924 15
rect -1947 -21 -1924 -15
rect -1868 15 -1845 21
rect -1868 -15 -1865 15
rect -1848 -15 -1845 15
rect -1868 -21 -1845 -15
rect -1789 15 -1766 21
rect -1789 -15 -1786 15
rect -1769 -15 -1766 15
rect -1789 -21 -1766 -15
rect -1710 15 -1687 21
rect -1710 -15 -1707 15
rect -1690 -15 -1687 15
rect -1710 -21 -1687 -15
rect -1631 15 -1608 21
rect -1631 -15 -1628 15
rect -1611 -15 -1608 15
rect -1631 -21 -1608 -15
rect -1552 15 -1529 21
rect -1552 -15 -1549 15
rect -1532 -15 -1529 15
rect -1552 -21 -1529 -15
rect -1473 15 -1450 21
rect -1473 -15 -1470 15
rect -1453 -15 -1450 15
rect -1473 -21 -1450 -15
rect -1394 15 -1371 21
rect -1394 -15 -1391 15
rect -1374 -15 -1371 15
rect -1394 -21 -1371 -15
rect -1315 15 -1292 21
rect -1315 -15 -1312 15
rect -1295 -15 -1292 15
rect -1315 -21 -1292 -15
rect -1236 15 -1213 21
rect -1236 -15 -1233 15
rect -1216 -15 -1213 15
rect -1236 -21 -1213 -15
rect -1157 15 -1134 21
rect -1157 -15 -1154 15
rect -1137 -15 -1134 15
rect -1157 -21 -1134 -15
rect -1078 15 -1055 21
rect -1078 -15 -1075 15
rect -1058 -15 -1055 15
rect -1078 -21 -1055 -15
rect -999 15 -976 21
rect -999 -15 -996 15
rect -979 -15 -976 15
rect -999 -21 -976 -15
rect -920 15 -897 21
rect -920 -15 -917 15
rect -900 -15 -897 15
rect -920 -21 -897 -15
rect -841 15 -818 21
rect -841 -15 -838 15
rect -821 -15 -818 15
rect -841 -21 -818 -15
rect -762 15 -739 21
rect -762 -15 -759 15
rect -742 -15 -739 15
rect -762 -21 -739 -15
rect -683 15 -660 21
rect -683 -15 -680 15
rect -663 -15 -660 15
rect -683 -21 -660 -15
rect -604 15 -581 21
rect -604 -15 -601 15
rect -584 -15 -581 15
rect -604 -21 -581 -15
rect -525 15 -502 21
rect -525 -15 -522 15
rect -505 -15 -502 15
rect -525 -21 -502 -15
rect -446 15 -423 21
rect -446 -15 -443 15
rect -426 -15 -423 15
rect -446 -21 -423 -15
rect -367 15 -344 21
rect -367 -15 -364 15
rect -347 -15 -344 15
rect -367 -21 -344 -15
rect -288 15 -265 21
rect -288 -15 -285 15
rect -268 -15 -265 15
rect -288 -21 -265 -15
rect -209 15 -186 21
rect -209 -15 -206 15
rect -189 -15 -186 15
rect -209 -21 -186 -15
rect -130 15 -107 21
rect -130 -15 -127 15
rect -110 -15 -107 15
rect -130 -21 -107 -15
rect -51 15 -28 21
rect -51 -15 -48 15
rect -31 -15 -28 15
rect -51 -21 -28 -15
rect 28 15 51 21
rect 28 -15 31 15
rect 48 -15 51 15
rect 28 -21 51 -15
rect 107 15 130 21
rect 107 -15 110 15
rect 127 -15 130 15
rect 107 -21 130 -15
rect 186 15 209 21
rect 186 -15 189 15
rect 206 -15 209 15
rect 186 -21 209 -15
rect 265 15 288 21
rect 265 -15 268 15
rect 285 -15 288 15
rect 265 -21 288 -15
rect 344 15 367 21
rect 344 -15 347 15
rect 364 -15 367 15
rect 344 -21 367 -15
rect 423 15 446 21
rect 423 -15 426 15
rect 443 -15 446 15
rect 423 -21 446 -15
rect 502 15 525 21
rect 502 -15 505 15
rect 522 -15 525 15
rect 502 -21 525 -15
rect 581 15 604 21
rect 581 -15 584 15
rect 601 -15 604 15
rect 581 -21 604 -15
rect 660 15 683 21
rect 660 -15 663 15
rect 680 -15 683 15
rect 660 -21 683 -15
rect 739 15 762 21
rect 739 -15 742 15
rect 759 -15 762 15
rect 739 -21 762 -15
rect 818 15 841 21
rect 818 -15 821 15
rect 838 -15 841 15
rect 818 -21 841 -15
rect 897 15 920 21
rect 897 -15 900 15
rect 917 -15 920 15
rect 897 -21 920 -15
rect 976 15 999 21
rect 976 -15 979 15
rect 996 -15 999 15
rect 976 -21 999 -15
rect 1055 15 1078 21
rect 1055 -15 1058 15
rect 1075 -15 1078 15
rect 1055 -21 1078 -15
rect 1134 15 1157 21
rect 1134 -15 1137 15
rect 1154 -15 1157 15
rect 1134 -21 1157 -15
rect 1213 15 1236 21
rect 1213 -15 1216 15
rect 1233 -15 1236 15
rect 1213 -21 1236 -15
rect 1292 15 1315 21
rect 1292 -15 1295 15
rect 1312 -15 1315 15
rect 1292 -21 1315 -15
rect 1371 15 1394 21
rect 1371 -15 1374 15
rect 1391 -15 1394 15
rect 1371 -21 1394 -15
rect 1450 15 1473 21
rect 1450 -15 1453 15
rect 1470 -15 1473 15
rect 1450 -21 1473 -15
rect 1529 15 1552 21
rect 1529 -15 1532 15
rect 1549 -15 1552 15
rect 1529 -21 1552 -15
rect 1608 15 1631 21
rect 1608 -15 1611 15
rect 1628 -15 1631 15
rect 1608 -21 1631 -15
rect 1687 15 1710 21
rect 1687 -15 1690 15
rect 1707 -15 1710 15
rect 1687 -21 1710 -15
rect 1766 15 1789 21
rect 1766 -15 1769 15
rect 1786 -15 1789 15
rect 1766 -21 1789 -15
rect 1845 15 1868 21
rect 1845 -15 1848 15
rect 1865 -15 1868 15
rect 1845 -21 1868 -15
rect 1924 15 1947 21
rect 1924 -15 1927 15
rect 1944 -15 1947 15
rect 1924 -21 1947 -15
rect 2003 15 2026 21
rect 2003 -15 2006 15
rect 2023 -15 2026 15
rect 2003 -21 2026 -15
rect -1998 -40 -1952 -37
rect -1998 -57 -1992 -40
rect -1958 -57 -1952 -40
rect -1998 -60 -1952 -57
rect -1919 -40 -1873 -37
rect -1919 -57 -1913 -40
rect -1879 -57 -1873 -40
rect -1919 -60 -1873 -57
rect -1840 -40 -1794 -37
rect -1840 -57 -1834 -40
rect -1800 -57 -1794 -40
rect -1840 -60 -1794 -57
rect -1761 -40 -1715 -37
rect -1761 -57 -1755 -40
rect -1721 -57 -1715 -40
rect -1761 -60 -1715 -57
rect -1682 -40 -1636 -37
rect -1682 -57 -1676 -40
rect -1642 -57 -1636 -40
rect -1682 -60 -1636 -57
rect -1603 -40 -1557 -37
rect -1603 -57 -1597 -40
rect -1563 -57 -1557 -40
rect -1603 -60 -1557 -57
rect -1524 -40 -1478 -37
rect -1524 -57 -1518 -40
rect -1484 -57 -1478 -40
rect -1524 -60 -1478 -57
rect -1445 -40 -1399 -37
rect -1445 -57 -1439 -40
rect -1405 -57 -1399 -40
rect -1445 -60 -1399 -57
rect -1366 -40 -1320 -37
rect -1366 -57 -1360 -40
rect -1326 -57 -1320 -40
rect -1366 -60 -1320 -57
rect -1287 -40 -1241 -37
rect -1287 -57 -1281 -40
rect -1247 -57 -1241 -40
rect -1287 -60 -1241 -57
rect -1208 -40 -1162 -37
rect -1208 -57 -1202 -40
rect -1168 -57 -1162 -40
rect -1208 -60 -1162 -57
rect -1129 -40 -1083 -37
rect -1129 -57 -1123 -40
rect -1089 -57 -1083 -40
rect -1129 -60 -1083 -57
rect -1050 -40 -1004 -37
rect -1050 -57 -1044 -40
rect -1010 -57 -1004 -40
rect -1050 -60 -1004 -57
rect -971 -40 -925 -37
rect -971 -57 -965 -40
rect -931 -57 -925 -40
rect -971 -60 -925 -57
rect -892 -40 -846 -37
rect -892 -57 -886 -40
rect -852 -57 -846 -40
rect -892 -60 -846 -57
rect -813 -40 -767 -37
rect -813 -57 -807 -40
rect -773 -57 -767 -40
rect -813 -60 -767 -57
rect -734 -40 -688 -37
rect -734 -57 -728 -40
rect -694 -57 -688 -40
rect -734 -60 -688 -57
rect -655 -40 -609 -37
rect -655 -57 -649 -40
rect -615 -57 -609 -40
rect -655 -60 -609 -57
rect -576 -40 -530 -37
rect -576 -57 -570 -40
rect -536 -57 -530 -40
rect -576 -60 -530 -57
rect -497 -40 -451 -37
rect -497 -57 -491 -40
rect -457 -57 -451 -40
rect -497 -60 -451 -57
rect -418 -40 -372 -37
rect -418 -57 -412 -40
rect -378 -57 -372 -40
rect -418 -60 -372 -57
rect -339 -40 -293 -37
rect -339 -57 -333 -40
rect -299 -57 -293 -40
rect -339 -60 -293 -57
rect -260 -40 -214 -37
rect -260 -57 -254 -40
rect -220 -57 -214 -40
rect -260 -60 -214 -57
rect -181 -40 -135 -37
rect -181 -57 -175 -40
rect -141 -57 -135 -40
rect -181 -60 -135 -57
rect -102 -40 -56 -37
rect -102 -57 -96 -40
rect -62 -57 -56 -40
rect -102 -60 -56 -57
rect -23 -40 23 -37
rect -23 -57 -17 -40
rect 17 -57 23 -40
rect -23 -60 23 -57
rect 56 -40 102 -37
rect 56 -57 62 -40
rect 96 -57 102 -40
rect 56 -60 102 -57
rect 135 -40 181 -37
rect 135 -57 141 -40
rect 175 -57 181 -40
rect 135 -60 181 -57
rect 214 -40 260 -37
rect 214 -57 220 -40
rect 254 -57 260 -40
rect 214 -60 260 -57
rect 293 -40 339 -37
rect 293 -57 299 -40
rect 333 -57 339 -40
rect 293 -60 339 -57
rect 372 -40 418 -37
rect 372 -57 378 -40
rect 412 -57 418 -40
rect 372 -60 418 -57
rect 451 -40 497 -37
rect 451 -57 457 -40
rect 491 -57 497 -40
rect 451 -60 497 -57
rect 530 -40 576 -37
rect 530 -57 536 -40
rect 570 -57 576 -40
rect 530 -60 576 -57
rect 609 -40 655 -37
rect 609 -57 615 -40
rect 649 -57 655 -40
rect 609 -60 655 -57
rect 688 -40 734 -37
rect 688 -57 694 -40
rect 728 -57 734 -40
rect 688 -60 734 -57
rect 767 -40 813 -37
rect 767 -57 773 -40
rect 807 -57 813 -40
rect 767 -60 813 -57
rect 846 -40 892 -37
rect 846 -57 852 -40
rect 886 -57 892 -40
rect 846 -60 892 -57
rect 925 -40 971 -37
rect 925 -57 931 -40
rect 965 -57 971 -40
rect 925 -60 971 -57
rect 1004 -40 1050 -37
rect 1004 -57 1010 -40
rect 1044 -57 1050 -40
rect 1004 -60 1050 -57
rect 1083 -40 1129 -37
rect 1083 -57 1089 -40
rect 1123 -57 1129 -40
rect 1083 -60 1129 -57
rect 1162 -40 1208 -37
rect 1162 -57 1168 -40
rect 1202 -57 1208 -40
rect 1162 -60 1208 -57
rect 1241 -40 1287 -37
rect 1241 -57 1247 -40
rect 1281 -57 1287 -40
rect 1241 -60 1287 -57
rect 1320 -40 1366 -37
rect 1320 -57 1326 -40
rect 1360 -57 1366 -40
rect 1320 -60 1366 -57
rect 1399 -40 1445 -37
rect 1399 -57 1405 -40
rect 1439 -57 1445 -40
rect 1399 -60 1445 -57
rect 1478 -40 1524 -37
rect 1478 -57 1484 -40
rect 1518 -57 1524 -40
rect 1478 -60 1524 -57
rect 1557 -40 1603 -37
rect 1557 -57 1563 -40
rect 1597 -57 1603 -40
rect 1557 -60 1603 -57
rect 1636 -40 1682 -37
rect 1636 -57 1642 -40
rect 1676 -57 1682 -40
rect 1636 -60 1682 -57
rect 1715 -40 1761 -37
rect 1715 -57 1721 -40
rect 1755 -57 1761 -40
rect 1715 -60 1761 -57
rect 1794 -40 1840 -37
rect 1794 -57 1800 -40
rect 1834 -57 1840 -40
rect 1794 -60 1840 -57
rect 1873 -40 1919 -37
rect 1873 -57 1879 -40
rect 1913 -57 1919 -40
rect 1873 -60 1919 -57
rect 1952 -40 1998 -37
rect 1952 -57 1958 -40
rect 1992 -57 1998 -40
rect 1952 -60 1998 -57
<< properties >>
string FIXED_BBOX -2081 -117 2081 117
string gencell sky130_fd_pr__nfet_03v3_nvt
string library sky130
string parameters w 0.42 l 0.5 m 1 nf 51 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
