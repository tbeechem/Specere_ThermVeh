magic
tech sky130A
magscale 1 2
timestamp 1717261150
<< error_s >>
rect 582 82 640 88
rect 582 48 594 82
rect 582 42 640 48
rect 582 -228 640 -222
rect 582 -262 594 -228
rect 582 -268 640 -262
<< metal1 >>
rect -600 -200 -400 0
rect 1600 -200 1800 0
rect 400 -1400 600 -1200
use sky130_fd_pr__nfet_01v8_648S5X  XM3
timestamp 1717261150
transform 1 0 611 0 1 -90
box -211 -310 211 310
<< labels >>
flabel metal1 1600 -200 1800 0 0 FreeSans 256 0 0 0 VLow_Src
port 2 nsew
flabel metal1 -600 -200 -400 0 0 FreeSans 256 0 0 0 VD_H
port 0 nsew
flabel metal1 400 -1400 600 -1200 0 FreeSans 256 0 0 0 VG_H
port 1 nsew
<< end >>
