magic
tech sky130A
magscale 1 2
timestamp 1717546687
<< metal1 >>
rect 5996 12654 7448 13018
rect 5996 11830 6392 12654
rect 7118 11830 7448 12654
rect 5996 6595 7448 11830
rect -7140 -2410 -6050 -135
rect 9920 -1540 10790 -385
rect -7140 -3506 -6050 -3500
rect -5260 -1925 -906 -1725
rect -5260 -6325 -5060 -1925
rect 9920 -2416 10790 -2410
rect -6088 -11910 -4636 -6325
rect -6088 -12734 -5758 -11910
rect -5032 -12734 -4636 -11910
rect -6088 -13328 -4636 -12734
<< via1 >>
rect 6392 11830 7118 12654
rect -7140 -3500 -6050 -2410
rect 9920 -2410 10790 -1540
rect -5758 -12734 -5032 -11910
<< metal2 >>
rect 6030 14670 7350 15100
rect 6030 13944 6392 14670
rect 7084 13944 7350 14670
rect 6030 12654 7350 13944
rect 6030 11830 6392 12654
rect 7118 11830 7350 12654
rect 6030 11468 7350 11830
rect -1290 7795 -305 7965
rect -1290 7050 -1120 7795
rect -440 7050 -305 7795
rect -1290 6370 -305 7050
rect 2430 7825 3430 7915
rect 2430 7080 2600 7825
rect 3280 7080 3430 7825
rect -965 4755 -765 6370
rect 2430 6320 3430 7080
rect 2805 4755 3005 6320
rect -965 4555 3005 4755
rect 1641 60 1841 4555
rect -8744 -3500 -8735 -2410
rect -7645 -3500 -7140 -2410
rect -6050 -3500 -6044 -2410
rect 1371 -2510 1581 -1795
rect 9914 -2410 9920 -1540
rect 10790 -2410 10796 -1540
rect -920 -2720 3040 -2510
rect -920 -5200 -710 -2720
rect 2830 -5175 3040 -2720
rect 9920 -2840 10790 -2410
rect 9920 -3719 10790 -3710
rect -1360 -7010 -325 -5200
rect -1360 -7755 -1205 -7010
rect -525 -7755 -325 -7010
rect 2395 -7010 3360 -5175
rect 2395 -7755 2565 -7010
rect 3245 -7755 3360 -7010
rect -1360 -7865 -325 -7755
rect -6054 -11910 -4734 -11742
rect -6054 -12734 -5758 -11910
rect -5032 -12734 -4734 -11910
rect -6054 -14352 -4734 -12734
rect -6054 -15078 -5790 -14352
rect -5098 -15078 -4734 -14352
rect -6054 -15374 -4734 -15078
<< via2 >>
rect 6392 13944 7084 14670
rect -1120 7050 -440 7795
rect 2600 7080 3280 7825
rect -8735 -3500 -7645 -2410
rect 9920 -3710 10790 -2840
rect -1205 -7755 -525 -7010
rect 2565 -7755 3245 -7010
rect -5790 -15078 -5098 -14352
<< metal3 >>
rect 6126 17284 7316 17692
rect 6126 16360 6352 17284
rect 7028 16360 7316 17284
rect 6126 14670 7316 16360
rect 6126 13944 6392 14670
rect 7084 13944 7316 14670
rect 6126 13596 7316 13944
rect -1260 9240 -300 9480
rect -1260 8460 -1080 9240
rect -420 8460 -300 9240
rect -1260 7795 -300 8460
rect -1260 7050 -1120 7795
rect -440 7050 -300 7795
rect -1260 6595 -300 7050
rect 2460 9240 3420 9480
rect 2460 8460 2640 9240
rect 3300 8460 3420 9240
rect 2460 7825 3420 8460
rect 2460 7080 2600 7825
rect 3280 7080 3420 7825
rect 2460 6595 3420 7080
rect -8740 -2410 -7640 -2405
rect -8740 -3500 -8735 -2410
rect -7645 -3500 -7640 -2410
rect -8740 -3505 -7640 -3500
rect 9915 -2840 10795 -2835
rect -8735 -4335 -7645 -3505
rect 9915 -3710 9920 -2840
rect 10790 -3710 10795 -2840
rect 9915 -3715 10795 -3710
rect -8735 -5431 -7645 -5425
rect 9920 -4730 10790 -3715
rect 9920 -5606 10790 -5600
rect -1325 -7010 -365 -6865
rect -1325 -7755 -1205 -7010
rect -525 -7475 -365 -7010
rect 2400 -7010 3360 -6920
rect -525 -7755 -360 -7475
rect -1325 -7825 -360 -7755
rect -1320 -9120 -360 -7825
rect -1320 -9900 -1140 -9120
rect -480 -9900 -360 -9120
rect -1320 -10140 -360 -9900
rect 2400 -7755 2565 -7010
rect 3245 -7755 3360 -7010
rect 2400 -9120 3360 -7755
rect 2400 -9900 2580 -9120
rect 3240 -9900 3360 -9120
rect 2400 -10140 3360 -9900
rect -6054 -14352 -4864 -14150
rect -6054 -15078 -5790 -14352
rect -5098 -15078 -4864 -14352
rect -6054 -17042 -4864 -15078
rect -6054 -17966 -5794 -17042
rect -5118 -17966 -4864 -17042
rect -6054 -18246 -4864 -17966
<< via3 >>
rect 6352 16360 7028 17284
rect -1080 8460 -420 9240
rect 2640 8460 3300 9240
rect -8735 -5425 -7645 -4335
rect 9920 -5600 10790 -4730
rect -1140 -9900 -480 -9120
rect 2580 -9900 3240 -9120
rect -5794 -17966 -5118 -17042
<< metal4 >>
rect 5418 24654 7998 25298
rect 5418 22976 5934 24654
rect 7354 22976 7998 24654
rect 5418 17284 7998 22976
rect 5418 16360 6352 17284
rect 7028 16360 7998 17284
rect 5418 15752 7998 16360
rect -1260 12660 -300 12900
rect -1260 12180 -1140 12660
rect -420 12180 -300 12660
rect -1260 9240 -300 12180
rect -1260 8460 -1080 9240
rect -420 8460 -300 9240
rect -1260 8100 -300 8460
rect 2460 12660 3420 12900
rect 2460 12180 2580 12660
rect 3300 12180 3420 12660
rect 2460 9240 3420 12180
rect 2460 8460 2640 9240
rect 3300 8460 3420 9240
rect 2460 8100 3420 8460
rect -8736 -4335 -7644 -4334
rect -8736 -5425 -8735 -4335
rect -7645 -5425 -7644 -4335
rect -8736 -5426 -7644 -5425
rect 9919 -4730 10791 -4729
rect -8735 -6240 -7645 -5426
rect 9919 -5600 9920 -4730
rect 10790 -5600 11785 -4730
rect 9919 -5601 10791 -5600
rect -1320 -9120 -360 -8760
rect -1320 -9900 -1140 -9120
rect -480 -9900 -360 -9120
rect -1320 -12840 -360 -9900
rect -1320 -13320 -1200 -12840
rect -480 -13320 -360 -12840
rect -1320 -13560 -360 -13320
rect 2400 -9120 3360 -8760
rect 2400 -9900 2580 -9120
rect 3240 -9900 3360 -9120
rect 2400 -12840 3360 -9900
rect 2400 -13320 2520 -12840
rect 3240 -13320 3360 -12840
rect 2400 -13560 3360 -13320
rect -6644 -17042 -4064 -16694
rect -6644 -17966 -5794 -17042
rect -5118 -17966 -4064 -17042
rect -6644 -23918 -4064 -17966
rect -6644 -25596 -6064 -23918
rect -4644 -25596 -4064 -23918
rect -6644 -26240 -4064 -25596
<< via4 >>
rect 5934 22976 7354 24654
rect -1140 12180 -420 12660
rect 2580 12180 3300 12660
rect 11785 -5600 12655 -4730
rect -8735 -7330 -7645 -6240
rect -1200 -13320 -480 -12840
rect 2520 -13320 3240 -12840
rect -6064 -25596 -4644 -23918
<< metal5 >>
rect -7104 25824 8896 42024
rect -28066 20160 -12066 25780
rect 5418 24654 7978 25824
rect 5418 22976 5934 24654
rect 7354 22976 7978 24654
rect 5418 22068 7978 22976
rect -28066 18900 -300 20160
rect 15120 20100 31120 25800
rect 14160 20084 31120 20100
rect 2392 18968 31120 20084
rect 2392 18952 5438 18968
rect 14160 18960 31120 18968
rect -28066 17000 -12066 18900
rect -28200 16000 -12060 17000
rect -28066 9580 -12066 16000
rect -1274 13080 -306 18900
rect -1294 12660 -284 13080
rect -1294 12180 -1140 12660
rect -420 12180 -284 12660
rect -1294 11980 -284 12180
rect 2426 12660 3436 18952
rect 2426 12180 2580 12660
rect 3300 12180 3436 12660
rect 2426 11980 3436 12180
rect 15120 9600 31120 18960
rect -28000 -86 -12000 7100
rect 15030 54 31030 7066
rect -28000 -1376 -11970 -86
rect -28000 -6240 -12000 -1376
rect 15015 -1486 31030 54
rect 11761 -4730 12679 -4706
rect 15030 -4730 31030 -1486
rect 11761 -5600 11785 -4730
rect 12655 -5600 31030 -4730
rect 11761 -5624 12679 -5600
rect -8759 -6240 -7621 -6216
rect -28000 -7330 -8735 -6240
rect -7645 -7330 -7621 -6240
rect -28000 -9100 -12000 -7330
rect -8759 -7354 -7621 -7330
rect 15030 -9134 31030 -5600
rect -28080 -19776 -12080 -11622
rect -1354 -12840 -344 -12640
rect -1354 -13320 -1200 -12840
rect -480 -13320 -344 -12840
rect -1354 -13740 -344 -13320
rect 2366 -12840 3376 -12640
rect 2366 -13320 2520 -12840
rect 3240 -13320 3376 -12840
rect -1334 -19776 -366 -13740
rect 2366 -19612 3376 -13320
rect 2332 -19628 5378 -19612
rect 15030 -19628 31030 -11764
rect -28080 -20702 -326 -19776
rect -28080 -27822 -12080 -20702
rect 2332 -20744 31030 -19628
rect 15002 -20852 31030 -20744
rect -6592 -23918 -4032 -23134
rect -6592 -25596 -6064 -23918
rect -4644 -25596 -4032 -23918
rect -6592 -27864 -4032 -25596
rect -7616 -44064 8384 -27864
rect 15030 -27964 31030 -20852
<< glass >>
rect -6800 26200 8600 41600
rect -27600 9800 -12466 25380
rect 15520 10000 30600 25400
rect -27600 -8700 -12400 6700
rect 15430 -8734 30630 6666
rect -27680 -27400 -12480 -12020
rect 15430 -27564 30630 -12164
rect -7200 -43800 8000 -28200
<< fillblock >>
rect -5298 -1240 9502 -240
use GSense_nFET_6Contacts_V2  GSense_nFET_3VD_3Vg_5nf_V2_0
timestamp 1717352107
transform 1 0 315 0 1 -138
box 0 0 1 1
use GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline  GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0
timestamp 1717386517
transform 1 0 -5224 0 1 -135
box -1366 -1870 15678 395
<< end >>
