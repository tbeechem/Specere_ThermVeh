magic
tech sky130A
timestamp 1717383051
<< pwell >>
rect -3589 -150 3589 150
<< nnmos >>
rect -3475 -21 -3425 21
rect -3337 -21 -3287 21
rect -3199 -21 -3149 21
rect -3061 -21 -3011 21
rect -2923 -21 -2873 21
rect -2785 -21 -2735 21
rect -2647 -21 -2597 21
rect -2509 -21 -2459 21
rect -2371 -21 -2321 21
rect -2233 -21 -2183 21
rect -2095 -21 -2045 21
rect -1957 -21 -1907 21
rect -1819 -21 -1769 21
rect -1681 -21 -1631 21
rect -1543 -21 -1493 21
rect -1405 -21 -1355 21
rect -1267 -21 -1217 21
rect -1129 -21 -1079 21
rect -991 -21 -941 21
rect -853 -21 -803 21
rect -715 -21 -665 21
rect -577 -21 -527 21
rect -439 -21 -389 21
rect -301 -21 -251 21
rect -163 -21 -113 21
rect -25 -21 25 21
rect 113 -21 163 21
rect 251 -21 301 21
rect 389 -21 439 21
rect 527 -21 577 21
rect 665 -21 715 21
rect 803 -21 853 21
rect 941 -21 991 21
rect 1079 -21 1129 21
rect 1217 -21 1267 21
rect 1355 -21 1405 21
rect 1493 -21 1543 21
rect 1631 -21 1681 21
rect 1769 -21 1819 21
rect 1907 -21 1957 21
rect 2045 -21 2095 21
rect 2183 -21 2233 21
rect 2321 -21 2371 21
rect 2459 -21 2509 21
rect 2597 -21 2647 21
rect 2735 -21 2785 21
rect 2873 -21 2923 21
rect 3011 -21 3061 21
rect 3149 -21 3199 21
rect 3287 -21 3337 21
rect 3425 -21 3475 21
<< mvndiff >>
rect -3504 15 -3475 21
rect -3504 -15 -3498 15
rect -3481 -15 -3475 15
rect -3504 -21 -3475 -15
rect -3425 15 -3396 21
rect -3425 -15 -3419 15
rect -3402 -15 -3396 15
rect -3425 -21 -3396 -15
rect -3366 15 -3337 21
rect -3366 -15 -3360 15
rect -3343 -15 -3337 15
rect -3366 -21 -3337 -15
rect -3287 15 -3258 21
rect -3287 -15 -3281 15
rect -3264 -15 -3258 15
rect -3287 -21 -3258 -15
rect -3228 15 -3199 21
rect -3228 -15 -3222 15
rect -3205 -15 -3199 15
rect -3228 -21 -3199 -15
rect -3149 15 -3120 21
rect -3149 -15 -3143 15
rect -3126 -15 -3120 15
rect -3149 -21 -3120 -15
rect -3090 15 -3061 21
rect -3090 -15 -3084 15
rect -3067 -15 -3061 15
rect -3090 -21 -3061 -15
rect -3011 15 -2982 21
rect -3011 -15 -3005 15
rect -2988 -15 -2982 15
rect -3011 -21 -2982 -15
rect -2952 15 -2923 21
rect -2952 -15 -2946 15
rect -2929 -15 -2923 15
rect -2952 -21 -2923 -15
rect -2873 15 -2844 21
rect -2873 -15 -2867 15
rect -2850 -15 -2844 15
rect -2873 -21 -2844 -15
rect -2814 15 -2785 21
rect -2814 -15 -2808 15
rect -2791 -15 -2785 15
rect -2814 -21 -2785 -15
rect -2735 15 -2706 21
rect -2735 -15 -2729 15
rect -2712 -15 -2706 15
rect -2735 -21 -2706 -15
rect -2676 15 -2647 21
rect -2676 -15 -2670 15
rect -2653 -15 -2647 15
rect -2676 -21 -2647 -15
rect -2597 15 -2568 21
rect -2597 -15 -2591 15
rect -2574 -15 -2568 15
rect -2597 -21 -2568 -15
rect -2538 15 -2509 21
rect -2538 -15 -2532 15
rect -2515 -15 -2509 15
rect -2538 -21 -2509 -15
rect -2459 15 -2430 21
rect -2459 -15 -2453 15
rect -2436 -15 -2430 15
rect -2459 -21 -2430 -15
rect -2400 15 -2371 21
rect -2400 -15 -2394 15
rect -2377 -15 -2371 15
rect -2400 -21 -2371 -15
rect -2321 15 -2292 21
rect -2321 -15 -2315 15
rect -2298 -15 -2292 15
rect -2321 -21 -2292 -15
rect -2262 15 -2233 21
rect -2262 -15 -2256 15
rect -2239 -15 -2233 15
rect -2262 -21 -2233 -15
rect -2183 15 -2154 21
rect -2183 -15 -2177 15
rect -2160 -15 -2154 15
rect -2183 -21 -2154 -15
rect -2124 15 -2095 21
rect -2124 -15 -2118 15
rect -2101 -15 -2095 15
rect -2124 -21 -2095 -15
rect -2045 15 -2016 21
rect -2045 -15 -2039 15
rect -2022 -15 -2016 15
rect -2045 -21 -2016 -15
rect -1986 15 -1957 21
rect -1986 -15 -1980 15
rect -1963 -15 -1957 15
rect -1986 -21 -1957 -15
rect -1907 15 -1878 21
rect -1907 -15 -1901 15
rect -1884 -15 -1878 15
rect -1907 -21 -1878 -15
rect -1848 15 -1819 21
rect -1848 -15 -1842 15
rect -1825 -15 -1819 15
rect -1848 -21 -1819 -15
rect -1769 15 -1740 21
rect -1769 -15 -1763 15
rect -1746 -15 -1740 15
rect -1769 -21 -1740 -15
rect -1710 15 -1681 21
rect -1710 -15 -1704 15
rect -1687 -15 -1681 15
rect -1710 -21 -1681 -15
rect -1631 15 -1602 21
rect -1631 -15 -1625 15
rect -1608 -15 -1602 15
rect -1631 -21 -1602 -15
rect -1572 15 -1543 21
rect -1572 -15 -1566 15
rect -1549 -15 -1543 15
rect -1572 -21 -1543 -15
rect -1493 15 -1464 21
rect -1493 -15 -1487 15
rect -1470 -15 -1464 15
rect -1493 -21 -1464 -15
rect -1434 15 -1405 21
rect -1434 -15 -1428 15
rect -1411 -15 -1405 15
rect -1434 -21 -1405 -15
rect -1355 15 -1326 21
rect -1355 -15 -1349 15
rect -1332 -15 -1326 15
rect -1355 -21 -1326 -15
rect -1296 15 -1267 21
rect -1296 -15 -1290 15
rect -1273 -15 -1267 15
rect -1296 -21 -1267 -15
rect -1217 15 -1188 21
rect -1217 -15 -1211 15
rect -1194 -15 -1188 15
rect -1217 -21 -1188 -15
rect -1158 15 -1129 21
rect -1158 -15 -1152 15
rect -1135 -15 -1129 15
rect -1158 -21 -1129 -15
rect -1079 15 -1050 21
rect -1079 -15 -1073 15
rect -1056 -15 -1050 15
rect -1079 -21 -1050 -15
rect -1020 15 -991 21
rect -1020 -15 -1014 15
rect -997 -15 -991 15
rect -1020 -21 -991 -15
rect -941 15 -912 21
rect -941 -15 -935 15
rect -918 -15 -912 15
rect -941 -21 -912 -15
rect -882 15 -853 21
rect -882 -15 -876 15
rect -859 -15 -853 15
rect -882 -21 -853 -15
rect -803 15 -774 21
rect -803 -15 -797 15
rect -780 -15 -774 15
rect -803 -21 -774 -15
rect -744 15 -715 21
rect -744 -15 -738 15
rect -721 -15 -715 15
rect -744 -21 -715 -15
rect -665 15 -636 21
rect -665 -15 -659 15
rect -642 -15 -636 15
rect -665 -21 -636 -15
rect -606 15 -577 21
rect -606 -15 -600 15
rect -583 -15 -577 15
rect -606 -21 -577 -15
rect -527 15 -498 21
rect -527 -15 -521 15
rect -504 -15 -498 15
rect -527 -21 -498 -15
rect -468 15 -439 21
rect -468 -15 -462 15
rect -445 -15 -439 15
rect -468 -21 -439 -15
rect -389 15 -360 21
rect -389 -15 -383 15
rect -366 -15 -360 15
rect -389 -21 -360 -15
rect -330 15 -301 21
rect -330 -15 -324 15
rect -307 -15 -301 15
rect -330 -21 -301 -15
rect -251 15 -222 21
rect -251 -15 -245 15
rect -228 -15 -222 15
rect -251 -21 -222 -15
rect -192 15 -163 21
rect -192 -15 -186 15
rect -169 -15 -163 15
rect -192 -21 -163 -15
rect -113 15 -84 21
rect -113 -15 -107 15
rect -90 -15 -84 15
rect -113 -21 -84 -15
rect -54 15 -25 21
rect -54 -15 -48 15
rect -31 -15 -25 15
rect -54 -21 -25 -15
rect 25 15 54 21
rect 25 -15 31 15
rect 48 -15 54 15
rect 25 -21 54 -15
rect 84 15 113 21
rect 84 -15 90 15
rect 107 -15 113 15
rect 84 -21 113 -15
rect 163 15 192 21
rect 163 -15 169 15
rect 186 -15 192 15
rect 163 -21 192 -15
rect 222 15 251 21
rect 222 -15 228 15
rect 245 -15 251 15
rect 222 -21 251 -15
rect 301 15 330 21
rect 301 -15 307 15
rect 324 -15 330 15
rect 301 -21 330 -15
rect 360 15 389 21
rect 360 -15 366 15
rect 383 -15 389 15
rect 360 -21 389 -15
rect 439 15 468 21
rect 439 -15 445 15
rect 462 -15 468 15
rect 439 -21 468 -15
rect 498 15 527 21
rect 498 -15 504 15
rect 521 -15 527 15
rect 498 -21 527 -15
rect 577 15 606 21
rect 577 -15 583 15
rect 600 -15 606 15
rect 577 -21 606 -15
rect 636 15 665 21
rect 636 -15 642 15
rect 659 -15 665 15
rect 636 -21 665 -15
rect 715 15 744 21
rect 715 -15 721 15
rect 738 -15 744 15
rect 715 -21 744 -15
rect 774 15 803 21
rect 774 -15 780 15
rect 797 -15 803 15
rect 774 -21 803 -15
rect 853 15 882 21
rect 853 -15 859 15
rect 876 -15 882 15
rect 853 -21 882 -15
rect 912 15 941 21
rect 912 -15 918 15
rect 935 -15 941 15
rect 912 -21 941 -15
rect 991 15 1020 21
rect 991 -15 997 15
rect 1014 -15 1020 15
rect 991 -21 1020 -15
rect 1050 15 1079 21
rect 1050 -15 1056 15
rect 1073 -15 1079 15
rect 1050 -21 1079 -15
rect 1129 15 1158 21
rect 1129 -15 1135 15
rect 1152 -15 1158 15
rect 1129 -21 1158 -15
rect 1188 15 1217 21
rect 1188 -15 1194 15
rect 1211 -15 1217 15
rect 1188 -21 1217 -15
rect 1267 15 1296 21
rect 1267 -15 1273 15
rect 1290 -15 1296 15
rect 1267 -21 1296 -15
rect 1326 15 1355 21
rect 1326 -15 1332 15
rect 1349 -15 1355 15
rect 1326 -21 1355 -15
rect 1405 15 1434 21
rect 1405 -15 1411 15
rect 1428 -15 1434 15
rect 1405 -21 1434 -15
rect 1464 15 1493 21
rect 1464 -15 1470 15
rect 1487 -15 1493 15
rect 1464 -21 1493 -15
rect 1543 15 1572 21
rect 1543 -15 1549 15
rect 1566 -15 1572 15
rect 1543 -21 1572 -15
rect 1602 15 1631 21
rect 1602 -15 1608 15
rect 1625 -15 1631 15
rect 1602 -21 1631 -15
rect 1681 15 1710 21
rect 1681 -15 1687 15
rect 1704 -15 1710 15
rect 1681 -21 1710 -15
rect 1740 15 1769 21
rect 1740 -15 1746 15
rect 1763 -15 1769 15
rect 1740 -21 1769 -15
rect 1819 15 1848 21
rect 1819 -15 1825 15
rect 1842 -15 1848 15
rect 1819 -21 1848 -15
rect 1878 15 1907 21
rect 1878 -15 1884 15
rect 1901 -15 1907 15
rect 1878 -21 1907 -15
rect 1957 15 1986 21
rect 1957 -15 1963 15
rect 1980 -15 1986 15
rect 1957 -21 1986 -15
rect 2016 15 2045 21
rect 2016 -15 2022 15
rect 2039 -15 2045 15
rect 2016 -21 2045 -15
rect 2095 15 2124 21
rect 2095 -15 2101 15
rect 2118 -15 2124 15
rect 2095 -21 2124 -15
rect 2154 15 2183 21
rect 2154 -15 2160 15
rect 2177 -15 2183 15
rect 2154 -21 2183 -15
rect 2233 15 2262 21
rect 2233 -15 2239 15
rect 2256 -15 2262 15
rect 2233 -21 2262 -15
rect 2292 15 2321 21
rect 2292 -15 2298 15
rect 2315 -15 2321 15
rect 2292 -21 2321 -15
rect 2371 15 2400 21
rect 2371 -15 2377 15
rect 2394 -15 2400 15
rect 2371 -21 2400 -15
rect 2430 15 2459 21
rect 2430 -15 2436 15
rect 2453 -15 2459 15
rect 2430 -21 2459 -15
rect 2509 15 2538 21
rect 2509 -15 2515 15
rect 2532 -15 2538 15
rect 2509 -21 2538 -15
rect 2568 15 2597 21
rect 2568 -15 2574 15
rect 2591 -15 2597 15
rect 2568 -21 2597 -15
rect 2647 15 2676 21
rect 2647 -15 2653 15
rect 2670 -15 2676 15
rect 2647 -21 2676 -15
rect 2706 15 2735 21
rect 2706 -15 2712 15
rect 2729 -15 2735 15
rect 2706 -21 2735 -15
rect 2785 15 2814 21
rect 2785 -15 2791 15
rect 2808 -15 2814 15
rect 2785 -21 2814 -15
rect 2844 15 2873 21
rect 2844 -15 2850 15
rect 2867 -15 2873 15
rect 2844 -21 2873 -15
rect 2923 15 2952 21
rect 2923 -15 2929 15
rect 2946 -15 2952 15
rect 2923 -21 2952 -15
rect 2982 15 3011 21
rect 2982 -15 2988 15
rect 3005 -15 3011 15
rect 2982 -21 3011 -15
rect 3061 15 3090 21
rect 3061 -15 3067 15
rect 3084 -15 3090 15
rect 3061 -21 3090 -15
rect 3120 15 3149 21
rect 3120 -15 3126 15
rect 3143 -15 3149 15
rect 3120 -21 3149 -15
rect 3199 15 3228 21
rect 3199 -15 3205 15
rect 3222 -15 3228 15
rect 3199 -21 3228 -15
rect 3258 15 3287 21
rect 3258 -15 3264 15
rect 3281 -15 3287 15
rect 3258 -21 3287 -15
rect 3337 15 3366 21
rect 3337 -15 3343 15
rect 3360 -15 3366 15
rect 3337 -21 3366 -15
rect 3396 15 3425 21
rect 3396 -15 3402 15
rect 3419 -15 3425 15
rect 3396 -21 3425 -15
rect 3475 15 3504 21
rect 3475 -15 3481 15
rect 3498 -15 3504 15
rect 3475 -21 3504 -15
<< mvndiffc >>
rect -3498 -15 -3481 15
rect -3419 -15 -3402 15
rect -3360 -15 -3343 15
rect -3281 -15 -3264 15
rect -3222 -15 -3205 15
rect -3143 -15 -3126 15
rect -3084 -15 -3067 15
rect -3005 -15 -2988 15
rect -2946 -15 -2929 15
rect -2867 -15 -2850 15
rect -2808 -15 -2791 15
rect -2729 -15 -2712 15
rect -2670 -15 -2653 15
rect -2591 -15 -2574 15
rect -2532 -15 -2515 15
rect -2453 -15 -2436 15
rect -2394 -15 -2377 15
rect -2315 -15 -2298 15
rect -2256 -15 -2239 15
rect -2177 -15 -2160 15
rect -2118 -15 -2101 15
rect -2039 -15 -2022 15
rect -1980 -15 -1963 15
rect -1901 -15 -1884 15
rect -1842 -15 -1825 15
rect -1763 -15 -1746 15
rect -1704 -15 -1687 15
rect -1625 -15 -1608 15
rect -1566 -15 -1549 15
rect -1487 -15 -1470 15
rect -1428 -15 -1411 15
rect -1349 -15 -1332 15
rect -1290 -15 -1273 15
rect -1211 -15 -1194 15
rect -1152 -15 -1135 15
rect -1073 -15 -1056 15
rect -1014 -15 -997 15
rect -935 -15 -918 15
rect -876 -15 -859 15
rect -797 -15 -780 15
rect -738 -15 -721 15
rect -659 -15 -642 15
rect -600 -15 -583 15
rect -521 -15 -504 15
rect -462 -15 -445 15
rect -383 -15 -366 15
rect -324 -15 -307 15
rect -245 -15 -228 15
rect -186 -15 -169 15
rect -107 -15 -90 15
rect -48 -15 -31 15
rect 31 -15 48 15
rect 90 -15 107 15
rect 169 -15 186 15
rect 228 -15 245 15
rect 307 -15 324 15
rect 366 -15 383 15
rect 445 -15 462 15
rect 504 -15 521 15
rect 583 -15 600 15
rect 642 -15 659 15
rect 721 -15 738 15
rect 780 -15 797 15
rect 859 -15 876 15
rect 918 -15 935 15
rect 997 -15 1014 15
rect 1056 -15 1073 15
rect 1135 -15 1152 15
rect 1194 -15 1211 15
rect 1273 -15 1290 15
rect 1332 -15 1349 15
rect 1411 -15 1428 15
rect 1470 -15 1487 15
rect 1549 -15 1566 15
rect 1608 -15 1625 15
rect 1687 -15 1704 15
rect 1746 -15 1763 15
rect 1825 -15 1842 15
rect 1884 -15 1901 15
rect 1963 -15 1980 15
rect 2022 -15 2039 15
rect 2101 -15 2118 15
rect 2160 -15 2177 15
rect 2239 -15 2256 15
rect 2298 -15 2315 15
rect 2377 -15 2394 15
rect 2436 -15 2453 15
rect 2515 -15 2532 15
rect 2574 -15 2591 15
rect 2653 -15 2670 15
rect 2712 -15 2729 15
rect 2791 -15 2808 15
rect 2850 -15 2867 15
rect 2929 -15 2946 15
rect 2988 -15 3005 15
rect 3067 -15 3084 15
rect 3126 -15 3143 15
rect 3205 -15 3222 15
rect 3264 -15 3281 15
rect 3343 -15 3360 15
rect 3402 -15 3419 15
rect 3481 -15 3498 15
<< mvpsubdiff >>
rect -3571 103 3571 132
rect -3571 -103 -3542 103
rect 3542 78 3571 103
rect 3542 -78 3548 78
rect 3565 -78 3571 78
rect 3542 -103 3571 -78
rect -3571 -132 3571 -103
<< mvpsubdiffcont >>
rect 3548 -78 3565 78
<< poly >>
rect -3475 57 -3425 65
rect -3475 40 -3467 57
rect -3433 40 -3425 57
rect -3475 21 -3425 40
rect -3337 57 -3287 65
rect -3337 40 -3329 57
rect -3295 40 -3287 57
rect -3337 21 -3287 40
rect -3199 57 -3149 65
rect -3199 40 -3191 57
rect -3157 40 -3149 57
rect -3199 21 -3149 40
rect -3061 57 -3011 65
rect -3061 40 -3053 57
rect -3019 40 -3011 57
rect -3061 21 -3011 40
rect -2923 57 -2873 65
rect -2923 40 -2915 57
rect -2881 40 -2873 57
rect -2923 21 -2873 40
rect -2785 57 -2735 65
rect -2785 40 -2777 57
rect -2743 40 -2735 57
rect -2785 21 -2735 40
rect -2647 57 -2597 65
rect -2647 40 -2639 57
rect -2605 40 -2597 57
rect -2647 21 -2597 40
rect -2509 57 -2459 65
rect -2509 40 -2501 57
rect -2467 40 -2459 57
rect -2509 21 -2459 40
rect -2371 57 -2321 65
rect -2371 40 -2363 57
rect -2329 40 -2321 57
rect -2371 21 -2321 40
rect -2233 57 -2183 65
rect -2233 40 -2225 57
rect -2191 40 -2183 57
rect -2233 21 -2183 40
rect -2095 57 -2045 65
rect -2095 40 -2087 57
rect -2053 40 -2045 57
rect -2095 21 -2045 40
rect -1957 57 -1907 65
rect -1957 40 -1949 57
rect -1915 40 -1907 57
rect -1957 21 -1907 40
rect -1819 57 -1769 65
rect -1819 40 -1811 57
rect -1777 40 -1769 57
rect -1819 21 -1769 40
rect -1681 57 -1631 65
rect -1681 40 -1673 57
rect -1639 40 -1631 57
rect -1681 21 -1631 40
rect -1543 57 -1493 65
rect -1543 40 -1535 57
rect -1501 40 -1493 57
rect -1543 21 -1493 40
rect -1405 57 -1355 65
rect -1405 40 -1397 57
rect -1363 40 -1355 57
rect -1405 21 -1355 40
rect -1267 57 -1217 65
rect -1267 40 -1259 57
rect -1225 40 -1217 57
rect -1267 21 -1217 40
rect -1129 57 -1079 65
rect -1129 40 -1121 57
rect -1087 40 -1079 57
rect -1129 21 -1079 40
rect -991 57 -941 65
rect -991 40 -983 57
rect -949 40 -941 57
rect -991 21 -941 40
rect -853 57 -803 65
rect -853 40 -845 57
rect -811 40 -803 57
rect -853 21 -803 40
rect -715 57 -665 65
rect -715 40 -707 57
rect -673 40 -665 57
rect -715 21 -665 40
rect -577 57 -527 65
rect -577 40 -569 57
rect -535 40 -527 57
rect -577 21 -527 40
rect -439 57 -389 65
rect -439 40 -431 57
rect -397 40 -389 57
rect -439 21 -389 40
rect -301 57 -251 65
rect -301 40 -293 57
rect -259 40 -251 57
rect -301 21 -251 40
rect -163 57 -113 65
rect -163 40 -155 57
rect -121 40 -113 57
rect -163 21 -113 40
rect -25 57 25 65
rect -25 40 -17 57
rect 17 40 25 57
rect -25 21 25 40
rect 113 57 163 65
rect 113 40 121 57
rect 155 40 163 57
rect 113 21 163 40
rect 251 57 301 65
rect 251 40 259 57
rect 293 40 301 57
rect 251 21 301 40
rect 389 57 439 65
rect 389 40 397 57
rect 431 40 439 57
rect 389 21 439 40
rect 527 57 577 65
rect 527 40 535 57
rect 569 40 577 57
rect 527 21 577 40
rect 665 57 715 65
rect 665 40 673 57
rect 707 40 715 57
rect 665 21 715 40
rect 803 57 853 65
rect 803 40 811 57
rect 845 40 853 57
rect 803 21 853 40
rect 941 57 991 65
rect 941 40 949 57
rect 983 40 991 57
rect 941 21 991 40
rect 1079 57 1129 65
rect 1079 40 1087 57
rect 1121 40 1129 57
rect 1079 21 1129 40
rect 1217 57 1267 65
rect 1217 40 1225 57
rect 1259 40 1267 57
rect 1217 21 1267 40
rect 1355 57 1405 65
rect 1355 40 1363 57
rect 1397 40 1405 57
rect 1355 21 1405 40
rect 1493 57 1543 65
rect 1493 40 1501 57
rect 1535 40 1543 57
rect 1493 21 1543 40
rect 1631 57 1681 65
rect 1631 40 1639 57
rect 1673 40 1681 57
rect 1631 21 1681 40
rect 1769 57 1819 65
rect 1769 40 1777 57
rect 1811 40 1819 57
rect 1769 21 1819 40
rect 1907 57 1957 65
rect 1907 40 1915 57
rect 1949 40 1957 57
rect 1907 21 1957 40
rect 2045 57 2095 65
rect 2045 40 2053 57
rect 2087 40 2095 57
rect 2045 21 2095 40
rect 2183 57 2233 65
rect 2183 40 2191 57
rect 2225 40 2233 57
rect 2183 21 2233 40
rect 2321 57 2371 65
rect 2321 40 2329 57
rect 2363 40 2371 57
rect 2321 21 2371 40
rect 2459 57 2509 65
rect 2459 40 2467 57
rect 2501 40 2509 57
rect 2459 21 2509 40
rect 2597 57 2647 65
rect 2597 40 2605 57
rect 2639 40 2647 57
rect 2597 21 2647 40
rect 2735 57 2785 65
rect 2735 40 2743 57
rect 2777 40 2785 57
rect 2735 21 2785 40
rect 2873 57 2923 65
rect 2873 40 2881 57
rect 2915 40 2923 57
rect 2873 21 2923 40
rect 3011 57 3061 65
rect 3011 40 3019 57
rect 3053 40 3061 57
rect 3011 21 3061 40
rect 3149 57 3199 65
rect 3149 40 3157 57
rect 3191 40 3199 57
rect 3149 21 3199 40
rect 3287 57 3337 65
rect 3287 40 3295 57
rect 3329 40 3337 57
rect 3287 21 3337 40
rect 3425 57 3475 65
rect 3425 40 3433 57
rect 3467 40 3475 57
rect 3425 21 3475 40
rect -3475 -40 -3425 -21
rect -3475 -57 -3467 -40
rect -3433 -57 -3425 -40
rect -3475 -65 -3425 -57
rect -3337 -40 -3287 -21
rect -3337 -57 -3329 -40
rect -3295 -57 -3287 -40
rect -3337 -65 -3287 -57
rect -3199 -40 -3149 -21
rect -3199 -57 -3191 -40
rect -3157 -57 -3149 -40
rect -3199 -65 -3149 -57
rect -3061 -40 -3011 -21
rect -3061 -57 -3053 -40
rect -3019 -57 -3011 -40
rect -3061 -65 -3011 -57
rect -2923 -40 -2873 -21
rect -2923 -57 -2915 -40
rect -2881 -57 -2873 -40
rect -2923 -65 -2873 -57
rect -2785 -40 -2735 -21
rect -2785 -57 -2777 -40
rect -2743 -57 -2735 -40
rect -2785 -65 -2735 -57
rect -2647 -40 -2597 -21
rect -2647 -57 -2639 -40
rect -2605 -57 -2597 -40
rect -2647 -65 -2597 -57
rect -2509 -40 -2459 -21
rect -2509 -57 -2501 -40
rect -2467 -57 -2459 -40
rect -2509 -65 -2459 -57
rect -2371 -40 -2321 -21
rect -2371 -57 -2363 -40
rect -2329 -57 -2321 -40
rect -2371 -65 -2321 -57
rect -2233 -40 -2183 -21
rect -2233 -57 -2225 -40
rect -2191 -57 -2183 -40
rect -2233 -65 -2183 -57
rect -2095 -40 -2045 -21
rect -2095 -57 -2087 -40
rect -2053 -57 -2045 -40
rect -2095 -65 -2045 -57
rect -1957 -40 -1907 -21
rect -1957 -57 -1949 -40
rect -1915 -57 -1907 -40
rect -1957 -65 -1907 -57
rect -1819 -40 -1769 -21
rect -1819 -57 -1811 -40
rect -1777 -57 -1769 -40
rect -1819 -65 -1769 -57
rect -1681 -40 -1631 -21
rect -1681 -57 -1673 -40
rect -1639 -57 -1631 -40
rect -1681 -65 -1631 -57
rect -1543 -40 -1493 -21
rect -1543 -57 -1535 -40
rect -1501 -57 -1493 -40
rect -1543 -65 -1493 -57
rect -1405 -40 -1355 -21
rect -1405 -57 -1397 -40
rect -1363 -57 -1355 -40
rect -1405 -65 -1355 -57
rect -1267 -40 -1217 -21
rect -1267 -57 -1259 -40
rect -1225 -57 -1217 -40
rect -1267 -65 -1217 -57
rect -1129 -40 -1079 -21
rect -1129 -57 -1121 -40
rect -1087 -57 -1079 -40
rect -1129 -65 -1079 -57
rect -991 -40 -941 -21
rect -991 -57 -983 -40
rect -949 -57 -941 -40
rect -991 -65 -941 -57
rect -853 -40 -803 -21
rect -853 -57 -845 -40
rect -811 -57 -803 -40
rect -853 -65 -803 -57
rect -715 -40 -665 -21
rect -715 -57 -707 -40
rect -673 -57 -665 -40
rect -715 -65 -665 -57
rect -577 -40 -527 -21
rect -577 -57 -569 -40
rect -535 -57 -527 -40
rect -577 -65 -527 -57
rect -439 -40 -389 -21
rect -439 -57 -431 -40
rect -397 -57 -389 -40
rect -439 -65 -389 -57
rect -301 -40 -251 -21
rect -301 -57 -293 -40
rect -259 -57 -251 -40
rect -301 -65 -251 -57
rect -163 -40 -113 -21
rect -163 -57 -155 -40
rect -121 -57 -113 -40
rect -163 -65 -113 -57
rect -25 -40 25 -21
rect -25 -57 -17 -40
rect 17 -57 25 -40
rect -25 -65 25 -57
rect 113 -40 163 -21
rect 113 -57 121 -40
rect 155 -57 163 -40
rect 113 -65 163 -57
rect 251 -40 301 -21
rect 251 -57 259 -40
rect 293 -57 301 -40
rect 251 -65 301 -57
rect 389 -40 439 -21
rect 389 -57 397 -40
rect 431 -57 439 -40
rect 389 -65 439 -57
rect 527 -40 577 -21
rect 527 -57 535 -40
rect 569 -57 577 -40
rect 527 -65 577 -57
rect 665 -40 715 -21
rect 665 -57 673 -40
rect 707 -57 715 -40
rect 665 -65 715 -57
rect 803 -40 853 -21
rect 803 -57 811 -40
rect 845 -57 853 -40
rect 803 -65 853 -57
rect 941 -40 991 -21
rect 941 -57 949 -40
rect 983 -57 991 -40
rect 941 -65 991 -57
rect 1079 -40 1129 -21
rect 1079 -57 1087 -40
rect 1121 -57 1129 -40
rect 1079 -65 1129 -57
rect 1217 -40 1267 -21
rect 1217 -57 1225 -40
rect 1259 -57 1267 -40
rect 1217 -65 1267 -57
rect 1355 -40 1405 -21
rect 1355 -57 1363 -40
rect 1397 -57 1405 -40
rect 1355 -65 1405 -57
rect 1493 -40 1543 -21
rect 1493 -57 1501 -40
rect 1535 -57 1543 -40
rect 1493 -65 1543 -57
rect 1631 -40 1681 -21
rect 1631 -57 1639 -40
rect 1673 -57 1681 -40
rect 1631 -65 1681 -57
rect 1769 -40 1819 -21
rect 1769 -57 1777 -40
rect 1811 -57 1819 -40
rect 1769 -65 1819 -57
rect 1907 -40 1957 -21
rect 1907 -57 1915 -40
rect 1949 -57 1957 -40
rect 1907 -65 1957 -57
rect 2045 -40 2095 -21
rect 2045 -57 2053 -40
rect 2087 -57 2095 -40
rect 2045 -65 2095 -57
rect 2183 -40 2233 -21
rect 2183 -57 2191 -40
rect 2225 -57 2233 -40
rect 2183 -65 2233 -57
rect 2321 -40 2371 -21
rect 2321 -57 2329 -40
rect 2363 -57 2371 -40
rect 2321 -65 2371 -57
rect 2459 -40 2509 -21
rect 2459 -57 2467 -40
rect 2501 -57 2509 -40
rect 2459 -65 2509 -57
rect 2597 -40 2647 -21
rect 2597 -57 2605 -40
rect 2639 -57 2647 -40
rect 2597 -65 2647 -57
rect 2735 -40 2785 -21
rect 2735 -57 2743 -40
rect 2777 -57 2785 -40
rect 2735 -65 2785 -57
rect 2873 -40 2923 -21
rect 2873 -57 2881 -40
rect 2915 -57 2923 -40
rect 2873 -65 2923 -57
rect 3011 -40 3061 -21
rect 3011 -57 3019 -40
rect 3053 -57 3061 -40
rect 3011 -65 3061 -57
rect 3149 -40 3199 -21
rect 3149 -57 3157 -40
rect 3191 -57 3199 -40
rect 3149 -65 3199 -57
rect 3287 -40 3337 -21
rect 3287 -57 3295 -40
rect 3329 -57 3337 -40
rect 3287 -65 3337 -57
rect 3425 -40 3475 -21
rect 3425 -57 3433 -40
rect 3467 -57 3475 -40
rect 3425 -65 3475 -57
<< polycont >>
rect -3467 40 -3433 57
rect -3329 40 -3295 57
rect -3191 40 -3157 57
rect -3053 40 -3019 57
rect -2915 40 -2881 57
rect -2777 40 -2743 57
rect -2639 40 -2605 57
rect -2501 40 -2467 57
rect -2363 40 -2329 57
rect -2225 40 -2191 57
rect -2087 40 -2053 57
rect -1949 40 -1915 57
rect -1811 40 -1777 57
rect -1673 40 -1639 57
rect -1535 40 -1501 57
rect -1397 40 -1363 57
rect -1259 40 -1225 57
rect -1121 40 -1087 57
rect -983 40 -949 57
rect -845 40 -811 57
rect -707 40 -673 57
rect -569 40 -535 57
rect -431 40 -397 57
rect -293 40 -259 57
rect -155 40 -121 57
rect -17 40 17 57
rect 121 40 155 57
rect 259 40 293 57
rect 397 40 431 57
rect 535 40 569 57
rect 673 40 707 57
rect 811 40 845 57
rect 949 40 983 57
rect 1087 40 1121 57
rect 1225 40 1259 57
rect 1363 40 1397 57
rect 1501 40 1535 57
rect 1639 40 1673 57
rect 1777 40 1811 57
rect 1915 40 1949 57
rect 2053 40 2087 57
rect 2191 40 2225 57
rect 2329 40 2363 57
rect 2467 40 2501 57
rect 2605 40 2639 57
rect 2743 40 2777 57
rect 2881 40 2915 57
rect 3019 40 3053 57
rect 3157 40 3191 57
rect 3295 40 3329 57
rect 3433 40 3467 57
rect -3467 -57 -3433 -40
rect -3329 -57 -3295 -40
rect -3191 -57 -3157 -40
rect -3053 -57 -3019 -40
rect -2915 -57 -2881 -40
rect -2777 -57 -2743 -40
rect -2639 -57 -2605 -40
rect -2501 -57 -2467 -40
rect -2363 -57 -2329 -40
rect -2225 -57 -2191 -40
rect -2087 -57 -2053 -40
rect -1949 -57 -1915 -40
rect -1811 -57 -1777 -40
rect -1673 -57 -1639 -40
rect -1535 -57 -1501 -40
rect -1397 -57 -1363 -40
rect -1259 -57 -1225 -40
rect -1121 -57 -1087 -40
rect -983 -57 -949 -40
rect -845 -57 -811 -40
rect -707 -57 -673 -40
rect -569 -57 -535 -40
rect -431 -57 -397 -40
rect -293 -57 -259 -40
rect -155 -57 -121 -40
rect -17 -57 17 -40
rect 121 -57 155 -40
rect 259 -57 293 -40
rect 397 -57 431 -40
rect 535 -57 569 -40
rect 673 -57 707 -40
rect 811 -57 845 -40
rect 949 -57 983 -40
rect 1087 -57 1121 -40
rect 1225 -57 1259 -40
rect 1363 -57 1397 -40
rect 1501 -57 1535 -40
rect 1639 -57 1673 -40
rect 1777 -57 1811 -40
rect 1915 -57 1949 -40
rect 2053 -57 2087 -40
rect 2191 -57 2225 -40
rect 2329 -57 2363 -40
rect 2467 -57 2501 -40
rect 2605 -57 2639 -40
rect 2743 -57 2777 -40
rect 2881 -57 2915 -40
rect 3019 -57 3053 -40
rect 3157 -57 3191 -40
rect 3295 -57 3329 -40
rect 3433 -57 3467 -40
<< locali >>
rect 3548 78 3565 86
rect -3475 40 -3467 57
rect -3433 40 -3425 57
rect -3337 40 -3329 57
rect -3295 40 -3287 57
rect -3199 40 -3191 57
rect -3157 40 -3149 57
rect -3061 40 -3053 57
rect -3019 40 -3011 57
rect -2923 40 -2915 57
rect -2881 40 -2873 57
rect -2785 40 -2777 57
rect -2743 40 -2735 57
rect -2647 40 -2639 57
rect -2605 40 -2597 57
rect -2509 40 -2501 57
rect -2467 40 -2459 57
rect -2371 40 -2363 57
rect -2329 40 -2321 57
rect -2233 40 -2225 57
rect -2191 40 -2183 57
rect -2095 40 -2087 57
rect -2053 40 -2045 57
rect -1957 40 -1949 57
rect -1915 40 -1907 57
rect -1819 40 -1811 57
rect -1777 40 -1769 57
rect -1681 40 -1673 57
rect -1639 40 -1631 57
rect -1543 40 -1535 57
rect -1501 40 -1493 57
rect -1405 40 -1397 57
rect -1363 40 -1355 57
rect -1267 40 -1259 57
rect -1225 40 -1217 57
rect -1129 40 -1121 57
rect -1087 40 -1079 57
rect -991 40 -983 57
rect -949 40 -941 57
rect -853 40 -845 57
rect -811 40 -803 57
rect -715 40 -707 57
rect -673 40 -665 57
rect -577 40 -569 57
rect -535 40 -527 57
rect -439 40 -431 57
rect -397 40 -389 57
rect -301 40 -293 57
rect -259 40 -251 57
rect -163 40 -155 57
rect -121 40 -113 57
rect -25 40 -17 57
rect 17 40 25 57
rect 113 40 121 57
rect 155 40 163 57
rect 251 40 259 57
rect 293 40 301 57
rect 389 40 397 57
rect 431 40 439 57
rect 527 40 535 57
rect 569 40 577 57
rect 665 40 673 57
rect 707 40 715 57
rect 803 40 811 57
rect 845 40 853 57
rect 941 40 949 57
rect 983 40 991 57
rect 1079 40 1087 57
rect 1121 40 1129 57
rect 1217 40 1225 57
rect 1259 40 1267 57
rect 1355 40 1363 57
rect 1397 40 1405 57
rect 1493 40 1501 57
rect 1535 40 1543 57
rect 1631 40 1639 57
rect 1673 40 1681 57
rect 1769 40 1777 57
rect 1811 40 1819 57
rect 1907 40 1915 57
rect 1949 40 1957 57
rect 2045 40 2053 57
rect 2087 40 2095 57
rect 2183 40 2191 57
rect 2225 40 2233 57
rect 2321 40 2329 57
rect 2363 40 2371 57
rect 2459 40 2467 57
rect 2501 40 2509 57
rect 2597 40 2605 57
rect 2639 40 2647 57
rect 2735 40 2743 57
rect 2777 40 2785 57
rect 2873 40 2881 57
rect 2915 40 2923 57
rect 3011 40 3019 57
rect 3053 40 3061 57
rect 3149 40 3157 57
rect 3191 40 3199 57
rect 3287 40 3295 57
rect 3329 40 3337 57
rect 3425 40 3433 57
rect 3467 40 3475 57
rect -3498 15 -3481 23
rect -3498 -23 -3481 -15
rect -3419 15 -3402 23
rect -3419 -23 -3402 -15
rect -3360 15 -3343 23
rect -3360 -23 -3343 -15
rect -3281 15 -3264 23
rect -3281 -23 -3264 -15
rect -3222 15 -3205 23
rect -3222 -23 -3205 -15
rect -3143 15 -3126 23
rect -3143 -23 -3126 -15
rect -3084 15 -3067 23
rect -3084 -23 -3067 -15
rect -3005 15 -2988 23
rect -3005 -23 -2988 -15
rect -2946 15 -2929 23
rect -2946 -23 -2929 -15
rect -2867 15 -2850 23
rect -2867 -23 -2850 -15
rect -2808 15 -2791 23
rect -2808 -23 -2791 -15
rect -2729 15 -2712 23
rect -2729 -23 -2712 -15
rect -2670 15 -2653 23
rect -2670 -23 -2653 -15
rect -2591 15 -2574 23
rect -2591 -23 -2574 -15
rect -2532 15 -2515 23
rect -2532 -23 -2515 -15
rect -2453 15 -2436 23
rect -2453 -23 -2436 -15
rect -2394 15 -2377 23
rect -2394 -23 -2377 -15
rect -2315 15 -2298 23
rect -2315 -23 -2298 -15
rect -2256 15 -2239 23
rect -2256 -23 -2239 -15
rect -2177 15 -2160 23
rect -2177 -23 -2160 -15
rect -2118 15 -2101 23
rect -2118 -23 -2101 -15
rect -2039 15 -2022 23
rect -2039 -23 -2022 -15
rect -1980 15 -1963 23
rect -1980 -23 -1963 -15
rect -1901 15 -1884 23
rect -1901 -23 -1884 -15
rect -1842 15 -1825 23
rect -1842 -23 -1825 -15
rect -1763 15 -1746 23
rect -1763 -23 -1746 -15
rect -1704 15 -1687 23
rect -1704 -23 -1687 -15
rect -1625 15 -1608 23
rect -1625 -23 -1608 -15
rect -1566 15 -1549 23
rect -1566 -23 -1549 -15
rect -1487 15 -1470 23
rect -1487 -23 -1470 -15
rect -1428 15 -1411 23
rect -1428 -23 -1411 -15
rect -1349 15 -1332 23
rect -1349 -23 -1332 -15
rect -1290 15 -1273 23
rect -1290 -23 -1273 -15
rect -1211 15 -1194 23
rect -1211 -23 -1194 -15
rect -1152 15 -1135 23
rect -1152 -23 -1135 -15
rect -1073 15 -1056 23
rect -1073 -23 -1056 -15
rect -1014 15 -997 23
rect -1014 -23 -997 -15
rect -935 15 -918 23
rect -935 -23 -918 -15
rect -876 15 -859 23
rect -876 -23 -859 -15
rect -797 15 -780 23
rect -797 -23 -780 -15
rect -738 15 -721 23
rect -738 -23 -721 -15
rect -659 15 -642 23
rect -659 -23 -642 -15
rect -600 15 -583 23
rect -600 -23 -583 -15
rect -521 15 -504 23
rect -521 -23 -504 -15
rect -462 15 -445 23
rect -462 -23 -445 -15
rect -383 15 -366 23
rect -383 -23 -366 -15
rect -324 15 -307 23
rect -324 -23 -307 -15
rect -245 15 -228 23
rect -245 -23 -228 -15
rect -186 15 -169 23
rect -186 -23 -169 -15
rect -107 15 -90 23
rect -107 -23 -90 -15
rect -48 15 -31 23
rect -48 -23 -31 -15
rect 31 15 48 23
rect 31 -23 48 -15
rect 90 15 107 23
rect 90 -23 107 -15
rect 169 15 186 23
rect 169 -23 186 -15
rect 228 15 245 23
rect 228 -23 245 -15
rect 307 15 324 23
rect 307 -23 324 -15
rect 366 15 383 23
rect 366 -23 383 -15
rect 445 15 462 23
rect 445 -23 462 -15
rect 504 15 521 23
rect 504 -23 521 -15
rect 583 15 600 23
rect 583 -23 600 -15
rect 642 15 659 23
rect 642 -23 659 -15
rect 721 15 738 23
rect 721 -23 738 -15
rect 780 15 797 23
rect 780 -23 797 -15
rect 859 15 876 23
rect 859 -23 876 -15
rect 918 15 935 23
rect 918 -23 935 -15
rect 997 15 1014 23
rect 997 -23 1014 -15
rect 1056 15 1073 23
rect 1056 -23 1073 -15
rect 1135 15 1152 23
rect 1135 -23 1152 -15
rect 1194 15 1211 23
rect 1194 -23 1211 -15
rect 1273 15 1290 23
rect 1273 -23 1290 -15
rect 1332 15 1349 23
rect 1332 -23 1349 -15
rect 1411 15 1428 23
rect 1411 -23 1428 -15
rect 1470 15 1487 23
rect 1470 -23 1487 -15
rect 1549 15 1566 23
rect 1549 -23 1566 -15
rect 1608 15 1625 23
rect 1608 -23 1625 -15
rect 1687 15 1704 23
rect 1687 -23 1704 -15
rect 1746 15 1763 23
rect 1746 -23 1763 -15
rect 1825 15 1842 23
rect 1825 -23 1842 -15
rect 1884 15 1901 23
rect 1884 -23 1901 -15
rect 1963 15 1980 23
rect 1963 -23 1980 -15
rect 2022 15 2039 23
rect 2022 -23 2039 -15
rect 2101 15 2118 23
rect 2101 -23 2118 -15
rect 2160 15 2177 23
rect 2160 -23 2177 -15
rect 2239 15 2256 23
rect 2239 -23 2256 -15
rect 2298 15 2315 23
rect 2298 -23 2315 -15
rect 2377 15 2394 23
rect 2377 -23 2394 -15
rect 2436 15 2453 23
rect 2436 -23 2453 -15
rect 2515 15 2532 23
rect 2515 -23 2532 -15
rect 2574 15 2591 23
rect 2574 -23 2591 -15
rect 2653 15 2670 23
rect 2653 -23 2670 -15
rect 2712 15 2729 23
rect 2712 -23 2729 -15
rect 2791 15 2808 23
rect 2791 -23 2808 -15
rect 2850 15 2867 23
rect 2850 -23 2867 -15
rect 2929 15 2946 23
rect 2929 -23 2946 -15
rect 2988 15 3005 23
rect 2988 -23 3005 -15
rect 3067 15 3084 23
rect 3067 -23 3084 -15
rect 3126 15 3143 23
rect 3126 -23 3143 -15
rect 3205 15 3222 23
rect 3205 -23 3222 -15
rect 3264 15 3281 23
rect 3264 -23 3281 -15
rect 3343 15 3360 23
rect 3343 -23 3360 -15
rect 3402 15 3419 23
rect 3402 -23 3419 -15
rect 3481 15 3498 23
rect 3481 -23 3498 -15
rect -3475 -57 -3467 -40
rect -3433 -57 -3425 -40
rect -3337 -57 -3329 -40
rect -3295 -57 -3287 -40
rect -3199 -57 -3191 -40
rect -3157 -57 -3149 -40
rect -3061 -57 -3053 -40
rect -3019 -57 -3011 -40
rect -2923 -57 -2915 -40
rect -2881 -57 -2873 -40
rect -2785 -57 -2777 -40
rect -2743 -57 -2735 -40
rect -2647 -57 -2639 -40
rect -2605 -57 -2597 -40
rect -2509 -57 -2501 -40
rect -2467 -57 -2459 -40
rect -2371 -57 -2363 -40
rect -2329 -57 -2321 -40
rect -2233 -57 -2225 -40
rect -2191 -57 -2183 -40
rect -2095 -57 -2087 -40
rect -2053 -57 -2045 -40
rect -1957 -57 -1949 -40
rect -1915 -57 -1907 -40
rect -1819 -57 -1811 -40
rect -1777 -57 -1769 -40
rect -1681 -57 -1673 -40
rect -1639 -57 -1631 -40
rect -1543 -57 -1535 -40
rect -1501 -57 -1493 -40
rect -1405 -57 -1397 -40
rect -1363 -57 -1355 -40
rect -1267 -57 -1259 -40
rect -1225 -57 -1217 -40
rect -1129 -57 -1121 -40
rect -1087 -57 -1079 -40
rect -991 -57 -983 -40
rect -949 -57 -941 -40
rect -853 -57 -845 -40
rect -811 -57 -803 -40
rect -715 -57 -707 -40
rect -673 -57 -665 -40
rect -577 -57 -569 -40
rect -535 -57 -527 -40
rect -439 -57 -431 -40
rect -397 -57 -389 -40
rect -301 -57 -293 -40
rect -259 -57 -251 -40
rect -163 -57 -155 -40
rect -121 -57 -113 -40
rect -25 -57 -17 -40
rect 17 -57 25 -40
rect 113 -57 121 -40
rect 155 -57 163 -40
rect 251 -57 259 -40
rect 293 -57 301 -40
rect 389 -57 397 -40
rect 431 -57 439 -40
rect 527 -57 535 -40
rect 569 -57 577 -40
rect 665 -57 673 -40
rect 707 -57 715 -40
rect 803 -57 811 -40
rect 845 -57 853 -40
rect 941 -57 949 -40
rect 983 -57 991 -40
rect 1079 -57 1087 -40
rect 1121 -57 1129 -40
rect 1217 -57 1225 -40
rect 1259 -57 1267 -40
rect 1355 -57 1363 -40
rect 1397 -57 1405 -40
rect 1493 -57 1501 -40
rect 1535 -57 1543 -40
rect 1631 -57 1639 -40
rect 1673 -57 1681 -40
rect 1769 -57 1777 -40
rect 1811 -57 1819 -40
rect 1907 -57 1915 -40
rect 1949 -57 1957 -40
rect 2045 -57 2053 -40
rect 2087 -57 2095 -40
rect 2183 -57 2191 -40
rect 2225 -57 2233 -40
rect 2321 -57 2329 -40
rect 2363 -57 2371 -40
rect 2459 -57 2467 -40
rect 2501 -57 2509 -40
rect 2597 -57 2605 -40
rect 2639 -57 2647 -40
rect 2735 -57 2743 -40
rect 2777 -57 2785 -40
rect 2873 -57 2881 -40
rect 2915 -57 2923 -40
rect 3011 -57 3019 -40
rect 3053 -57 3061 -40
rect 3149 -57 3157 -40
rect 3191 -57 3199 -40
rect 3287 -57 3295 -40
rect 3329 -57 3337 -40
rect 3425 -57 3433 -40
rect 3467 -57 3475 -40
rect 3548 -86 3565 -78
<< viali >>
rect -3467 40 -3433 57
rect -3329 40 -3295 57
rect -3191 40 -3157 57
rect -3053 40 -3019 57
rect -2915 40 -2881 57
rect -2777 40 -2743 57
rect -2639 40 -2605 57
rect -2501 40 -2467 57
rect -2363 40 -2329 57
rect -2225 40 -2191 57
rect -2087 40 -2053 57
rect -1949 40 -1915 57
rect -1811 40 -1777 57
rect -1673 40 -1639 57
rect -1535 40 -1501 57
rect -1397 40 -1363 57
rect -1259 40 -1225 57
rect -1121 40 -1087 57
rect -983 40 -949 57
rect -845 40 -811 57
rect -707 40 -673 57
rect -569 40 -535 57
rect -431 40 -397 57
rect -293 40 -259 57
rect -155 40 -121 57
rect -17 40 17 57
rect 121 40 155 57
rect 259 40 293 57
rect 397 40 431 57
rect 535 40 569 57
rect 673 40 707 57
rect 811 40 845 57
rect 949 40 983 57
rect 1087 40 1121 57
rect 1225 40 1259 57
rect 1363 40 1397 57
rect 1501 40 1535 57
rect 1639 40 1673 57
rect 1777 40 1811 57
rect 1915 40 1949 57
rect 2053 40 2087 57
rect 2191 40 2225 57
rect 2329 40 2363 57
rect 2467 40 2501 57
rect 2605 40 2639 57
rect 2743 40 2777 57
rect 2881 40 2915 57
rect 3019 40 3053 57
rect 3157 40 3191 57
rect 3295 40 3329 57
rect 3433 40 3467 57
rect -3498 -15 -3481 15
rect -3419 -15 -3402 15
rect -3360 -15 -3343 15
rect -3281 -15 -3264 15
rect -3222 -15 -3205 15
rect -3143 -15 -3126 15
rect -3084 -15 -3067 15
rect -3005 -15 -2988 15
rect -2946 -15 -2929 15
rect -2867 -15 -2850 15
rect -2808 -15 -2791 15
rect -2729 -15 -2712 15
rect -2670 -15 -2653 15
rect -2591 -15 -2574 15
rect -2532 -15 -2515 15
rect -2453 -15 -2436 15
rect -2394 -15 -2377 15
rect -2315 -15 -2298 15
rect -2256 -15 -2239 15
rect -2177 -15 -2160 15
rect -2118 -15 -2101 15
rect -2039 -15 -2022 15
rect -1980 -15 -1963 15
rect -1901 -15 -1884 15
rect -1842 -15 -1825 15
rect -1763 -15 -1746 15
rect -1704 -15 -1687 15
rect -1625 -15 -1608 15
rect -1566 -15 -1549 15
rect -1487 -15 -1470 15
rect -1428 -15 -1411 15
rect -1349 -15 -1332 15
rect -1290 -15 -1273 15
rect -1211 -15 -1194 15
rect -1152 -15 -1135 15
rect -1073 -15 -1056 15
rect -1014 -15 -997 15
rect -935 -15 -918 15
rect -876 -15 -859 15
rect -797 -15 -780 15
rect -738 -15 -721 15
rect -659 -15 -642 15
rect -600 -15 -583 15
rect -521 -15 -504 15
rect -462 -15 -445 15
rect -383 -15 -366 15
rect -324 -15 -307 15
rect -245 -15 -228 15
rect -186 -15 -169 15
rect -107 -15 -90 15
rect -48 -15 -31 15
rect 31 -15 48 15
rect 90 -15 107 15
rect 169 -15 186 15
rect 228 -15 245 15
rect 307 -15 324 15
rect 366 -15 383 15
rect 445 -15 462 15
rect 504 -15 521 15
rect 583 -15 600 15
rect 642 -15 659 15
rect 721 -15 738 15
rect 780 -15 797 15
rect 859 -15 876 15
rect 918 -15 935 15
rect 997 -15 1014 15
rect 1056 -15 1073 15
rect 1135 -15 1152 15
rect 1194 -15 1211 15
rect 1273 -15 1290 15
rect 1332 -15 1349 15
rect 1411 -15 1428 15
rect 1470 -15 1487 15
rect 1549 -15 1566 15
rect 1608 -15 1625 15
rect 1687 -15 1704 15
rect 1746 -15 1763 15
rect 1825 -15 1842 15
rect 1884 -15 1901 15
rect 1963 -15 1980 15
rect 2022 -15 2039 15
rect 2101 -15 2118 15
rect 2160 -15 2177 15
rect 2239 -15 2256 15
rect 2298 -15 2315 15
rect 2377 -15 2394 15
rect 2436 -15 2453 15
rect 2515 -15 2532 15
rect 2574 -15 2591 15
rect 2653 -15 2670 15
rect 2712 -15 2729 15
rect 2791 -15 2808 15
rect 2850 -15 2867 15
rect 2929 -15 2946 15
rect 2988 -15 3005 15
rect 3067 -15 3084 15
rect 3126 -15 3143 15
rect 3205 -15 3222 15
rect 3264 -15 3281 15
rect 3343 -15 3360 15
rect 3402 -15 3419 15
rect 3481 -15 3498 15
rect -3467 -57 -3433 -40
rect -3329 -57 -3295 -40
rect -3191 -57 -3157 -40
rect -3053 -57 -3019 -40
rect -2915 -57 -2881 -40
rect -2777 -57 -2743 -40
rect -2639 -57 -2605 -40
rect -2501 -57 -2467 -40
rect -2363 -57 -2329 -40
rect -2225 -57 -2191 -40
rect -2087 -57 -2053 -40
rect -1949 -57 -1915 -40
rect -1811 -57 -1777 -40
rect -1673 -57 -1639 -40
rect -1535 -57 -1501 -40
rect -1397 -57 -1363 -40
rect -1259 -57 -1225 -40
rect -1121 -57 -1087 -40
rect -983 -57 -949 -40
rect -845 -57 -811 -40
rect -707 -57 -673 -40
rect -569 -57 -535 -40
rect -431 -57 -397 -40
rect -293 -57 -259 -40
rect -155 -57 -121 -40
rect -17 -57 17 -40
rect 121 -57 155 -40
rect 259 -57 293 -40
rect 397 -57 431 -40
rect 535 -57 569 -40
rect 673 -57 707 -40
rect 811 -57 845 -40
rect 949 -57 983 -40
rect 1087 -57 1121 -40
rect 1225 -57 1259 -40
rect 1363 -57 1397 -40
rect 1501 -57 1535 -40
rect 1639 -57 1673 -40
rect 1777 -57 1811 -40
rect 1915 -57 1949 -40
rect 2053 -57 2087 -40
rect 2191 -57 2225 -40
rect 2329 -57 2363 -40
rect 2467 -57 2501 -40
rect 2605 -57 2639 -40
rect 2743 -57 2777 -40
rect 2881 -57 2915 -40
rect 3019 -57 3053 -40
rect 3157 -57 3191 -40
rect 3295 -57 3329 -40
rect 3433 -57 3467 -40
<< metal1 >>
rect -3473 57 -3427 60
rect -3473 40 -3467 57
rect -3433 40 -3427 57
rect -3473 37 -3427 40
rect -3335 57 -3289 60
rect -3335 40 -3329 57
rect -3295 40 -3289 57
rect -3335 37 -3289 40
rect -3197 57 -3151 60
rect -3197 40 -3191 57
rect -3157 40 -3151 57
rect -3197 37 -3151 40
rect -3059 57 -3013 60
rect -3059 40 -3053 57
rect -3019 40 -3013 57
rect -3059 37 -3013 40
rect -2921 57 -2875 60
rect -2921 40 -2915 57
rect -2881 40 -2875 57
rect -2921 37 -2875 40
rect -2783 57 -2737 60
rect -2783 40 -2777 57
rect -2743 40 -2737 57
rect -2783 37 -2737 40
rect -2645 57 -2599 60
rect -2645 40 -2639 57
rect -2605 40 -2599 57
rect -2645 37 -2599 40
rect -2507 57 -2461 60
rect -2507 40 -2501 57
rect -2467 40 -2461 57
rect -2507 37 -2461 40
rect -2369 57 -2323 60
rect -2369 40 -2363 57
rect -2329 40 -2323 57
rect -2369 37 -2323 40
rect -2231 57 -2185 60
rect -2231 40 -2225 57
rect -2191 40 -2185 57
rect -2231 37 -2185 40
rect -2093 57 -2047 60
rect -2093 40 -2087 57
rect -2053 40 -2047 57
rect -2093 37 -2047 40
rect -1955 57 -1909 60
rect -1955 40 -1949 57
rect -1915 40 -1909 57
rect -1955 37 -1909 40
rect -1817 57 -1771 60
rect -1817 40 -1811 57
rect -1777 40 -1771 57
rect -1817 37 -1771 40
rect -1679 57 -1633 60
rect -1679 40 -1673 57
rect -1639 40 -1633 57
rect -1679 37 -1633 40
rect -1541 57 -1495 60
rect -1541 40 -1535 57
rect -1501 40 -1495 57
rect -1541 37 -1495 40
rect -1403 57 -1357 60
rect -1403 40 -1397 57
rect -1363 40 -1357 57
rect -1403 37 -1357 40
rect -1265 57 -1219 60
rect -1265 40 -1259 57
rect -1225 40 -1219 57
rect -1265 37 -1219 40
rect -1127 57 -1081 60
rect -1127 40 -1121 57
rect -1087 40 -1081 57
rect -1127 37 -1081 40
rect -989 57 -943 60
rect -989 40 -983 57
rect -949 40 -943 57
rect -989 37 -943 40
rect -851 57 -805 60
rect -851 40 -845 57
rect -811 40 -805 57
rect -851 37 -805 40
rect -713 57 -667 60
rect -713 40 -707 57
rect -673 40 -667 57
rect -713 37 -667 40
rect -575 57 -529 60
rect -575 40 -569 57
rect -535 40 -529 57
rect -575 37 -529 40
rect -437 57 -391 60
rect -437 40 -431 57
rect -397 40 -391 57
rect -437 37 -391 40
rect -299 57 -253 60
rect -299 40 -293 57
rect -259 40 -253 57
rect -299 37 -253 40
rect -161 57 -115 60
rect -161 40 -155 57
rect -121 40 -115 57
rect -161 37 -115 40
rect -23 57 23 60
rect -23 40 -17 57
rect 17 40 23 57
rect -23 37 23 40
rect 115 57 161 60
rect 115 40 121 57
rect 155 40 161 57
rect 115 37 161 40
rect 253 57 299 60
rect 253 40 259 57
rect 293 40 299 57
rect 253 37 299 40
rect 391 57 437 60
rect 391 40 397 57
rect 431 40 437 57
rect 391 37 437 40
rect 529 57 575 60
rect 529 40 535 57
rect 569 40 575 57
rect 529 37 575 40
rect 667 57 713 60
rect 667 40 673 57
rect 707 40 713 57
rect 667 37 713 40
rect 805 57 851 60
rect 805 40 811 57
rect 845 40 851 57
rect 805 37 851 40
rect 943 57 989 60
rect 943 40 949 57
rect 983 40 989 57
rect 943 37 989 40
rect 1081 57 1127 60
rect 1081 40 1087 57
rect 1121 40 1127 57
rect 1081 37 1127 40
rect 1219 57 1265 60
rect 1219 40 1225 57
rect 1259 40 1265 57
rect 1219 37 1265 40
rect 1357 57 1403 60
rect 1357 40 1363 57
rect 1397 40 1403 57
rect 1357 37 1403 40
rect 1495 57 1541 60
rect 1495 40 1501 57
rect 1535 40 1541 57
rect 1495 37 1541 40
rect 1633 57 1679 60
rect 1633 40 1639 57
rect 1673 40 1679 57
rect 1633 37 1679 40
rect 1771 57 1817 60
rect 1771 40 1777 57
rect 1811 40 1817 57
rect 1771 37 1817 40
rect 1909 57 1955 60
rect 1909 40 1915 57
rect 1949 40 1955 57
rect 1909 37 1955 40
rect 2047 57 2093 60
rect 2047 40 2053 57
rect 2087 40 2093 57
rect 2047 37 2093 40
rect 2185 57 2231 60
rect 2185 40 2191 57
rect 2225 40 2231 57
rect 2185 37 2231 40
rect 2323 57 2369 60
rect 2323 40 2329 57
rect 2363 40 2369 57
rect 2323 37 2369 40
rect 2461 57 2507 60
rect 2461 40 2467 57
rect 2501 40 2507 57
rect 2461 37 2507 40
rect 2599 57 2645 60
rect 2599 40 2605 57
rect 2639 40 2645 57
rect 2599 37 2645 40
rect 2737 57 2783 60
rect 2737 40 2743 57
rect 2777 40 2783 57
rect 2737 37 2783 40
rect 2875 57 2921 60
rect 2875 40 2881 57
rect 2915 40 2921 57
rect 2875 37 2921 40
rect 3013 57 3059 60
rect 3013 40 3019 57
rect 3053 40 3059 57
rect 3013 37 3059 40
rect 3151 57 3197 60
rect 3151 40 3157 57
rect 3191 40 3197 57
rect 3151 37 3197 40
rect 3289 57 3335 60
rect 3289 40 3295 57
rect 3329 40 3335 57
rect 3289 37 3335 40
rect 3427 57 3473 60
rect 3427 40 3433 57
rect 3467 40 3473 57
rect 3427 37 3473 40
rect -3501 15 -3478 21
rect -3501 -15 -3498 15
rect -3481 -15 -3478 15
rect -3501 -21 -3478 -15
rect -3422 15 -3399 21
rect -3422 -15 -3419 15
rect -3402 -15 -3399 15
rect -3422 -21 -3399 -15
rect -3363 15 -3340 21
rect -3363 -15 -3360 15
rect -3343 -15 -3340 15
rect -3363 -21 -3340 -15
rect -3284 15 -3261 21
rect -3284 -15 -3281 15
rect -3264 -15 -3261 15
rect -3284 -21 -3261 -15
rect -3225 15 -3202 21
rect -3225 -15 -3222 15
rect -3205 -15 -3202 15
rect -3225 -21 -3202 -15
rect -3146 15 -3123 21
rect -3146 -15 -3143 15
rect -3126 -15 -3123 15
rect -3146 -21 -3123 -15
rect -3087 15 -3064 21
rect -3087 -15 -3084 15
rect -3067 -15 -3064 15
rect -3087 -21 -3064 -15
rect -3008 15 -2985 21
rect -3008 -15 -3005 15
rect -2988 -15 -2985 15
rect -3008 -21 -2985 -15
rect -2949 15 -2926 21
rect -2949 -15 -2946 15
rect -2929 -15 -2926 15
rect -2949 -21 -2926 -15
rect -2870 15 -2847 21
rect -2870 -15 -2867 15
rect -2850 -15 -2847 15
rect -2870 -21 -2847 -15
rect -2811 15 -2788 21
rect -2811 -15 -2808 15
rect -2791 -15 -2788 15
rect -2811 -21 -2788 -15
rect -2732 15 -2709 21
rect -2732 -15 -2729 15
rect -2712 -15 -2709 15
rect -2732 -21 -2709 -15
rect -2673 15 -2650 21
rect -2673 -15 -2670 15
rect -2653 -15 -2650 15
rect -2673 -21 -2650 -15
rect -2594 15 -2571 21
rect -2594 -15 -2591 15
rect -2574 -15 -2571 15
rect -2594 -21 -2571 -15
rect -2535 15 -2512 21
rect -2535 -15 -2532 15
rect -2515 -15 -2512 15
rect -2535 -21 -2512 -15
rect -2456 15 -2433 21
rect -2456 -15 -2453 15
rect -2436 -15 -2433 15
rect -2456 -21 -2433 -15
rect -2397 15 -2374 21
rect -2397 -15 -2394 15
rect -2377 -15 -2374 15
rect -2397 -21 -2374 -15
rect -2318 15 -2295 21
rect -2318 -15 -2315 15
rect -2298 -15 -2295 15
rect -2318 -21 -2295 -15
rect -2259 15 -2236 21
rect -2259 -15 -2256 15
rect -2239 -15 -2236 15
rect -2259 -21 -2236 -15
rect -2180 15 -2157 21
rect -2180 -15 -2177 15
rect -2160 -15 -2157 15
rect -2180 -21 -2157 -15
rect -2121 15 -2098 21
rect -2121 -15 -2118 15
rect -2101 -15 -2098 15
rect -2121 -21 -2098 -15
rect -2042 15 -2019 21
rect -2042 -15 -2039 15
rect -2022 -15 -2019 15
rect -2042 -21 -2019 -15
rect -1983 15 -1960 21
rect -1983 -15 -1980 15
rect -1963 -15 -1960 15
rect -1983 -21 -1960 -15
rect -1904 15 -1881 21
rect -1904 -15 -1901 15
rect -1884 -15 -1881 15
rect -1904 -21 -1881 -15
rect -1845 15 -1822 21
rect -1845 -15 -1842 15
rect -1825 -15 -1822 15
rect -1845 -21 -1822 -15
rect -1766 15 -1743 21
rect -1766 -15 -1763 15
rect -1746 -15 -1743 15
rect -1766 -21 -1743 -15
rect -1707 15 -1684 21
rect -1707 -15 -1704 15
rect -1687 -15 -1684 15
rect -1707 -21 -1684 -15
rect -1628 15 -1605 21
rect -1628 -15 -1625 15
rect -1608 -15 -1605 15
rect -1628 -21 -1605 -15
rect -1569 15 -1546 21
rect -1569 -15 -1566 15
rect -1549 -15 -1546 15
rect -1569 -21 -1546 -15
rect -1490 15 -1467 21
rect -1490 -15 -1487 15
rect -1470 -15 -1467 15
rect -1490 -21 -1467 -15
rect -1431 15 -1408 21
rect -1431 -15 -1428 15
rect -1411 -15 -1408 15
rect -1431 -21 -1408 -15
rect -1352 15 -1329 21
rect -1352 -15 -1349 15
rect -1332 -15 -1329 15
rect -1352 -21 -1329 -15
rect -1293 15 -1270 21
rect -1293 -15 -1290 15
rect -1273 -15 -1270 15
rect -1293 -21 -1270 -15
rect -1214 15 -1191 21
rect -1214 -15 -1211 15
rect -1194 -15 -1191 15
rect -1214 -21 -1191 -15
rect -1155 15 -1132 21
rect -1155 -15 -1152 15
rect -1135 -15 -1132 15
rect -1155 -21 -1132 -15
rect -1076 15 -1053 21
rect -1076 -15 -1073 15
rect -1056 -15 -1053 15
rect -1076 -21 -1053 -15
rect -1017 15 -994 21
rect -1017 -15 -1014 15
rect -997 -15 -994 15
rect -1017 -21 -994 -15
rect -938 15 -915 21
rect -938 -15 -935 15
rect -918 -15 -915 15
rect -938 -21 -915 -15
rect -879 15 -856 21
rect -879 -15 -876 15
rect -859 -15 -856 15
rect -879 -21 -856 -15
rect -800 15 -777 21
rect -800 -15 -797 15
rect -780 -15 -777 15
rect -800 -21 -777 -15
rect -741 15 -718 21
rect -741 -15 -738 15
rect -721 -15 -718 15
rect -741 -21 -718 -15
rect -662 15 -639 21
rect -662 -15 -659 15
rect -642 -15 -639 15
rect -662 -21 -639 -15
rect -603 15 -580 21
rect -603 -15 -600 15
rect -583 -15 -580 15
rect -603 -21 -580 -15
rect -524 15 -501 21
rect -524 -15 -521 15
rect -504 -15 -501 15
rect -524 -21 -501 -15
rect -465 15 -442 21
rect -465 -15 -462 15
rect -445 -15 -442 15
rect -465 -21 -442 -15
rect -386 15 -363 21
rect -386 -15 -383 15
rect -366 -15 -363 15
rect -386 -21 -363 -15
rect -327 15 -304 21
rect -327 -15 -324 15
rect -307 -15 -304 15
rect -327 -21 -304 -15
rect -248 15 -225 21
rect -248 -15 -245 15
rect -228 -15 -225 15
rect -248 -21 -225 -15
rect -189 15 -166 21
rect -189 -15 -186 15
rect -169 -15 -166 15
rect -189 -21 -166 -15
rect -110 15 -87 21
rect -110 -15 -107 15
rect -90 -15 -87 15
rect -110 -21 -87 -15
rect -51 15 -28 21
rect -51 -15 -48 15
rect -31 -15 -28 15
rect -51 -21 -28 -15
rect 28 15 51 21
rect 28 -15 31 15
rect 48 -15 51 15
rect 28 -21 51 -15
rect 87 15 110 21
rect 87 -15 90 15
rect 107 -15 110 15
rect 87 -21 110 -15
rect 166 15 189 21
rect 166 -15 169 15
rect 186 -15 189 15
rect 166 -21 189 -15
rect 225 15 248 21
rect 225 -15 228 15
rect 245 -15 248 15
rect 225 -21 248 -15
rect 304 15 327 21
rect 304 -15 307 15
rect 324 -15 327 15
rect 304 -21 327 -15
rect 363 15 386 21
rect 363 -15 366 15
rect 383 -15 386 15
rect 363 -21 386 -15
rect 442 15 465 21
rect 442 -15 445 15
rect 462 -15 465 15
rect 442 -21 465 -15
rect 501 15 524 21
rect 501 -15 504 15
rect 521 -15 524 15
rect 501 -21 524 -15
rect 580 15 603 21
rect 580 -15 583 15
rect 600 -15 603 15
rect 580 -21 603 -15
rect 639 15 662 21
rect 639 -15 642 15
rect 659 -15 662 15
rect 639 -21 662 -15
rect 718 15 741 21
rect 718 -15 721 15
rect 738 -15 741 15
rect 718 -21 741 -15
rect 777 15 800 21
rect 777 -15 780 15
rect 797 -15 800 15
rect 777 -21 800 -15
rect 856 15 879 21
rect 856 -15 859 15
rect 876 -15 879 15
rect 856 -21 879 -15
rect 915 15 938 21
rect 915 -15 918 15
rect 935 -15 938 15
rect 915 -21 938 -15
rect 994 15 1017 21
rect 994 -15 997 15
rect 1014 -15 1017 15
rect 994 -21 1017 -15
rect 1053 15 1076 21
rect 1053 -15 1056 15
rect 1073 -15 1076 15
rect 1053 -21 1076 -15
rect 1132 15 1155 21
rect 1132 -15 1135 15
rect 1152 -15 1155 15
rect 1132 -21 1155 -15
rect 1191 15 1214 21
rect 1191 -15 1194 15
rect 1211 -15 1214 15
rect 1191 -21 1214 -15
rect 1270 15 1293 21
rect 1270 -15 1273 15
rect 1290 -15 1293 15
rect 1270 -21 1293 -15
rect 1329 15 1352 21
rect 1329 -15 1332 15
rect 1349 -15 1352 15
rect 1329 -21 1352 -15
rect 1408 15 1431 21
rect 1408 -15 1411 15
rect 1428 -15 1431 15
rect 1408 -21 1431 -15
rect 1467 15 1490 21
rect 1467 -15 1470 15
rect 1487 -15 1490 15
rect 1467 -21 1490 -15
rect 1546 15 1569 21
rect 1546 -15 1549 15
rect 1566 -15 1569 15
rect 1546 -21 1569 -15
rect 1605 15 1628 21
rect 1605 -15 1608 15
rect 1625 -15 1628 15
rect 1605 -21 1628 -15
rect 1684 15 1707 21
rect 1684 -15 1687 15
rect 1704 -15 1707 15
rect 1684 -21 1707 -15
rect 1743 15 1766 21
rect 1743 -15 1746 15
rect 1763 -15 1766 15
rect 1743 -21 1766 -15
rect 1822 15 1845 21
rect 1822 -15 1825 15
rect 1842 -15 1845 15
rect 1822 -21 1845 -15
rect 1881 15 1904 21
rect 1881 -15 1884 15
rect 1901 -15 1904 15
rect 1881 -21 1904 -15
rect 1960 15 1983 21
rect 1960 -15 1963 15
rect 1980 -15 1983 15
rect 1960 -21 1983 -15
rect 2019 15 2042 21
rect 2019 -15 2022 15
rect 2039 -15 2042 15
rect 2019 -21 2042 -15
rect 2098 15 2121 21
rect 2098 -15 2101 15
rect 2118 -15 2121 15
rect 2098 -21 2121 -15
rect 2157 15 2180 21
rect 2157 -15 2160 15
rect 2177 -15 2180 15
rect 2157 -21 2180 -15
rect 2236 15 2259 21
rect 2236 -15 2239 15
rect 2256 -15 2259 15
rect 2236 -21 2259 -15
rect 2295 15 2318 21
rect 2295 -15 2298 15
rect 2315 -15 2318 15
rect 2295 -21 2318 -15
rect 2374 15 2397 21
rect 2374 -15 2377 15
rect 2394 -15 2397 15
rect 2374 -21 2397 -15
rect 2433 15 2456 21
rect 2433 -15 2436 15
rect 2453 -15 2456 15
rect 2433 -21 2456 -15
rect 2512 15 2535 21
rect 2512 -15 2515 15
rect 2532 -15 2535 15
rect 2512 -21 2535 -15
rect 2571 15 2594 21
rect 2571 -15 2574 15
rect 2591 -15 2594 15
rect 2571 -21 2594 -15
rect 2650 15 2673 21
rect 2650 -15 2653 15
rect 2670 -15 2673 15
rect 2650 -21 2673 -15
rect 2709 15 2732 21
rect 2709 -15 2712 15
rect 2729 -15 2732 15
rect 2709 -21 2732 -15
rect 2788 15 2811 21
rect 2788 -15 2791 15
rect 2808 -15 2811 15
rect 2788 -21 2811 -15
rect 2847 15 2870 21
rect 2847 -15 2850 15
rect 2867 -15 2870 15
rect 2847 -21 2870 -15
rect 2926 15 2949 21
rect 2926 -15 2929 15
rect 2946 -15 2949 15
rect 2926 -21 2949 -15
rect 2985 15 3008 21
rect 2985 -15 2988 15
rect 3005 -15 3008 15
rect 2985 -21 3008 -15
rect 3064 15 3087 21
rect 3064 -15 3067 15
rect 3084 -15 3087 15
rect 3064 -21 3087 -15
rect 3123 15 3146 21
rect 3123 -15 3126 15
rect 3143 -15 3146 15
rect 3123 -21 3146 -15
rect 3202 15 3225 21
rect 3202 -15 3205 15
rect 3222 -15 3225 15
rect 3202 -21 3225 -15
rect 3261 15 3284 21
rect 3261 -15 3264 15
rect 3281 -15 3284 15
rect 3261 -21 3284 -15
rect 3340 15 3363 21
rect 3340 -15 3343 15
rect 3360 -15 3363 15
rect 3340 -21 3363 -15
rect 3399 15 3422 21
rect 3399 -15 3402 15
rect 3419 -15 3422 15
rect 3399 -21 3422 -15
rect 3478 15 3501 21
rect 3478 -15 3481 15
rect 3498 -15 3501 15
rect 3478 -21 3501 -15
rect -3473 -40 -3427 -37
rect -3473 -57 -3467 -40
rect -3433 -57 -3427 -40
rect -3473 -60 -3427 -57
rect -3335 -40 -3289 -37
rect -3335 -57 -3329 -40
rect -3295 -57 -3289 -40
rect -3335 -60 -3289 -57
rect -3197 -40 -3151 -37
rect -3197 -57 -3191 -40
rect -3157 -57 -3151 -40
rect -3197 -60 -3151 -57
rect -3059 -40 -3013 -37
rect -3059 -57 -3053 -40
rect -3019 -57 -3013 -40
rect -3059 -60 -3013 -57
rect -2921 -40 -2875 -37
rect -2921 -57 -2915 -40
rect -2881 -57 -2875 -40
rect -2921 -60 -2875 -57
rect -2783 -40 -2737 -37
rect -2783 -57 -2777 -40
rect -2743 -57 -2737 -40
rect -2783 -60 -2737 -57
rect -2645 -40 -2599 -37
rect -2645 -57 -2639 -40
rect -2605 -57 -2599 -40
rect -2645 -60 -2599 -57
rect -2507 -40 -2461 -37
rect -2507 -57 -2501 -40
rect -2467 -57 -2461 -40
rect -2507 -60 -2461 -57
rect -2369 -40 -2323 -37
rect -2369 -57 -2363 -40
rect -2329 -57 -2323 -40
rect -2369 -60 -2323 -57
rect -2231 -40 -2185 -37
rect -2231 -57 -2225 -40
rect -2191 -57 -2185 -40
rect -2231 -60 -2185 -57
rect -2093 -40 -2047 -37
rect -2093 -57 -2087 -40
rect -2053 -57 -2047 -40
rect -2093 -60 -2047 -57
rect -1955 -40 -1909 -37
rect -1955 -57 -1949 -40
rect -1915 -57 -1909 -40
rect -1955 -60 -1909 -57
rect -1817 -40 -1771 -37
rect -1817 -57 -1811 -40
rect -1777 -57 -1771 -40
rect -1817 -60 -1771 -57
rect -1679 -40 -1633 -37
rect -1679 -57 -1673 -40
rect -1639 -57 -1633 -40
rect -1679 -60 -1633 -57
rect -1541 -40 -1495 -37
rect -1541 -57 -1535 -40
rect -1501 -57 -1495 -40
rect -1541 -60 -1495 -57
rect -1403 -40 -1357 -37
rect -1403 -57 -1397 -40
rect -1363 -57 -1357 -40
rect -1403 -60 -1357 -57
rect -1265 -40 -1219 -37
rect -1265 -57 -1259 -40
rect -1225 -57 -1219 -40
rect -1265 -60 -1219 -57
rect -1127 -40 -1081 -37
rect -1127 -57 -1121 -40
rect -1087 -57 -1081 -40
rect -1127 -60 -1081 -57
rect -989 -40 -943 -37
rect -989 -57 -983 -40
rect -949 -57 -943 -40
rect -989 -60 -943 -57
rect -851 -40 -805 -37
rect -851 -57 -845 -40
rect -811 -57 -805 -40
rect -851 -60 -805 -57
rect -713 -40 -667 -37
rect -713 -57 -707 -40
rect -673 -57 -667 -40
rect -713 -60 -667 -57
rect -575 -40 -529 -37
rect -575 -57 -569 -40
rect -535 -57 -529 -40
rect -575 -60 -529 -57
rect -437 -40 -391 -37
rect -437 -57 -431 -40
rect -397 -57 -391 -40
rect -437 -60 -391 -57
rect -299 -40 -253 -37
rect -299 -57 -293 -40
rect -259 -57 -253 -40
rect -299 -60 -253 -57
rect -161 -40 -115 -37
rect -161 -57 -155 -40
rect -121 -57 -115 -40
rect -161 -60 -115 -57
rect -23 -40 23 -37
rect -23 -57 -17 -40
rect 17 -57 23 -40
rect -23 -60 23 -57
rect 115 -40 161 -37
rect 115 -57 121 -40
rect 155 -57 161 -40
rect 115 -60 161 -57
rect 253 -40 299 -37
rect 253 -57 259 -40
rect 293 -57 299 -40
rect 253 -60 299 -57
rect 391 -40 437 -37
rect 391 -57 397 -40
rect 431 -57 437 -40
rect 391 -60 437 -57
rect 529 -40 575 -37
rect 529 -57 535 -40
rect 569 -57 575 -40
rect 529 -60 575 -57
rect 667 -40 713 -37
rect 667 -57 673 -40
rect 707 -57 713 -40
rect 667 -60 713 -57
rect 805 -40 851 -37
rect 805 -57 811 -40
rect 845 -57 851 -40
rect 805 -60 851 -57
rect 943 -40 989 -37
rect 943 -57 949 -40
rect 983 -57 989 -40
rect 943 -60 989 -57
rect 1081 -40 1127 -37
rect 1081 -57 1087 -40
rect 1121 -57 1127 -40
rect 1081 -60 1127 -57
rect 1219 -40 1265 -37
rect 1219 -57 1225 -40
rect 1259 -57 1265 -40
rect 1219 -60 1265 -57
rect 1357 -40 1403 -37
rect 1357 -57 1363 -40
rect 1397 -57 1403 -40
rect 1357 -60 1403 -57
rect 1495 -40 1541 -37
rect 1495 -57 1501 -40
rect 1535 -57 1541 -40
rect 1495 -60 1541 -57
rect 1633 -40 1679 -37
rect 1633 -57 1639 -40
rect 1673 -57 1679 -40
rect 1633 -60 1679 -57
rect 1771 -40 1817 -37
rect 1771 -57 1777 -40
rect 1811 -57 1817 -40
rect 1771 -60 1817 -57
rect 1909 -40 1955 -37
rect 1909 -57 1915 -40
rect 1949 -57 1955 -40
rect 1909 -60 1955 -57
rect 2047 -40 2093 -37
rect 2047 -57 2053 -40
rect 2087 -57 2093 -40
rect 2047 -60 2093 -57
rect 2185 -40 2231 -37
rect 2185 -57 2191 -40
rect 2225 -57 2231 -40
rect 2185 -60 2231 -57
rect 2323 -40 2369 -37
rect 2323 -57 2329 -40
rect 2363 -57 2369 -40
rect 2323 -60 2369 -57
rect 2461 -40 2507 -37
rect 2461 -57 2467 -40
rect 2501 -57 2507 -40
rect 2461 -60 2507 -57
rect 2599 -40 2645 -37
rect 2599 -57 2605 -40
rect 2639 -57 2645 -40
rect 2599 -60 2645 -57
rect 2737 -40 2783 -37
rect 2737 -57 2743 -40
rect 2777 -57 2783 -40
rect 2737 -60 2783 -57
rect 2875 -40 2921 -37
rect 2875 -57 2881 -40
rect 2915 -57 2921 -40
rect 2875 -60 2921 -57
rect 3013 -40 3059 -37
rect 3013 -57 3019 -40
rect 3053 -57 3059 -40
rect 3013 -60 3059 -57
rect 3151 -40 3197 -37
rect 3151 -57 3157 -40
rect 3191 -57 3197 -40
rect 3151 -60 3197 -57
rect 3289 -40 3335 -37
rect 3289 -57 3295 -40
rect 3329 -57 3335 -40
rect 3289 -60 3335 -57
rect 3427 -40 3473 -37
rect 3427 -57 3433 -40
rect 3467 -57 3473 -40
rect 3427 -60 3473 -57
rect -3494 -124 -3406 -103
<< properties >>
string FIXED_BBOX -3556 -117 3556 117
string gencell sky130_fd_pr__nfet_03v3_nvt
string library sky130
string parameters w 0.42 l 0.5 m 1 nf 51 diffcov 100 polycov 100 guard 1 glc 0 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
