magic
tech sky130A
timestamp 1717352107
<< end >>
