magic
tech sky130A
magscale 1 2
timestamp 1717299026
<< error_p >>
rect 1980 -80 1986 -74
rect 2134 -80 2140 -74
rect 1974 -86 1980 -80
rect 2140 -86 2146 -80
rect 1974 -240 1980 -234
rect 2140 -240 2146 -234
rect 1980 -246 1986 -240
rect 2134 -246 2140 -240
<< metal1 >>
rect -1260 3260 -300 3420
rect -1260 2660 -1100 3260
rect -500 2660 -300 3260
rect -1260 1740 -300 2660
rect 2460 3260 3420 3420
rect 2460 2660 2620 3260
rect 3220 2660 3420 3260
rect 2460 1740 3420 2660
rect -1260 1140 3420 1740
rect -280 -80 160 -40
rect -280 -240 -220 -80
rect -60 -240 160 -80
rect -280 -280 160 -240
rect -1320 -2400 3360 -1800
rect -1320 -3320 -360 -2400
rect -1320 -3920 -1160 -3320
rect -560 -3920 -360 -3320
rect -1320 -4080 -360 -3920
rect 2400 -3320 3360 -2400
rect 2400 -3920 2560 -3320
rect 3160 -3920 3360 -3320
rect 2400 -4080 3360 -3920
<< via1 >>
rect -1100 2660 -500 3260
rect 2620 2660 3220 3260
rect -220 -240 -60 -80
rect 1980 -240 2140 -80
rect -1160 -3920 -560 -3320
rect 2560 -3920 3160 -3320
<< metal2 >>
rect -1260 6240 -300 6360
rect -1260 5580 -1080 6240
rect -420 5580 -300 6240
rect -1260 3260 -300 5580
rect -1260 2660 -1100 3260
rect -500 2660 -300 3260
rect 2460 6240 3420 6360
rect 2460 5580 2640 6240
rect 3300 5580 3420 6240
rect 2460 3260 3420 5580
rect 2460 2660 2620 3260
rect 3220 2660 3420 3260
rect -240 -80 -40 -60
rect -240 -240 -220 -80
rect -60 -240 -40 -80
rect -240 -840 -40 -240
rect 1960 -80 2160 -60
rect 1960 -240 1980 -80
rect 2140 -100 2160 -80
rect 2140 -110 2240 -100
rect 2140 -210 2690 -110
rect 2140 -220 2240 -210
rect 2140 -240 2160 -220
rect 1960 -260 2160 -240
rect 2590 -230 2690 -210
rect 3240 -200 3440 -180
rect 3240 -230 3260 -200
rect 2590 -330 3260 -230
rect 3240 -360 3260 -330
rect 3420 -360 3440 -200
rect 3240 -380 3440 -360
rect -880 -880 -40 -840
rect -880 -1000 -840 -880
rect -640 -1000 -40 -880
rect -880 -1040 -40 -1000
rect -1320 -3920 -1160 -3320
rect -560 -3920 -360 -3320
rect -1320 -6240 -360 -3920
rect -1320 -6900 -1140 -6240
rect -480 -6900 -360 -6240
rect -1320 -7020 -360 -6900
rect 2400 -3920 2560 -3320
rect 3160 -3920 3360 -3320
rect 2400 -6240 3360 -3920
rect 2400 -6900 2580 -6240
rect 3240 -6900 3360 -6240
rect 2400 -7020 3360 -6900
<< via2 >>
rect -1080 5580 -420 6240
rect 2640 5580 3300 6240
rect 3260 -360 3420 -200
rect -840 -1000 -640 -880
rect -1140 -6900 -480 -6240
rect 2580 -6900 3240 -6240
<< metal3 >>
rect -1260 9240 -300 9480
rect -1260 8460 -1080 9240
rect -420 8460 -300 9240
rect -1260 6240 -300 8460
rect -1260 5580 -1080 6240
rect -420 5580 -300 6240
rect -1260 5400 -300 5580
rect 2460 9240 3420 9480
rect 2460 8460 2640 9240
rect 3300 8460 3420 9240
rect 2460 6240 3420 8460
rect 2460 5580 2640 6240
rect 3300 5580 3420 6240
rect 2460 5400 3420 5580
rect -2564 -840 -1332 -82
rect 3240 -200 3460 -180
rect 3240 -360 3260 -200
rect 3420 -202 3460 -200
rect 3420 -319 4577 -202
rect 5373 -319 6247 -299
rect 3420 -356 6247 -319
rect 3420 -360 3460 -356
rect 3240 -380 3460 -360
rect 4423 -600 6247 -356
rect -2564 -1040 -2514 -840
rect -2314 -880 -600 -840
rect -2314 -1000 -840 -880
rect -640 -1000 -600 -880
rect 4423 -885 5550 -600
rect -2314 -1040 -600 -1000
rect -2564 -1390 -1332 -1040
rect 4419 -1050 5550 -885
rect 6000 -1050 6247 -600
rect 4419 -1335 6247 -1050
rect -1320 -6240 -360 -6060
rect -1320 -6900 -1140 -6240
rect -480 -6900 -360 -6240
rect -1320 -9120 -360 -6900
rect -1320 -9900 -1140 -9120
rect -480 -9900 -360 -9120
rect -1320 -10140 -360 -9900
rect 2400 -6240 3360 -6060
rect 2400 -6900 2580 -6240
rect 3240 -6900 3360 -6240
rect 2400 -9120 3360 -6900
rect 2400 -9900 2580 -9120
rect 3240 -9900 3360 -9120
rect 2400 -10140 3360 -9900
<< via3 >>
rect -1080 8460 -420 9240
rect 2640 8460 3300 9240
rect -2514 -1040 -2314 -840
rect 5550 -1050 6000 -600
rect -1140 -9900 -480 -9120
rect 2580 -9900 3240 -9120
<< metal4 >>
rect -1260 12660 -300 12900
rect -1260 12180 -1140 12660
rect -420 12180 -300 12660
rect -1260 9240 -300 12180
rect -1260 8460 -1080 9240
rect -420 8460 -300 9240
rect -1260 8100 -300 8460
rect 2460 12660 3420 12900
rect 2460 12180 2580 12660
rect 3300 12180 3420 12660
rect 2460 9240 3420 12180
rect 2460 8460 2640 9240
rect 3300 8460 3420 9240
rect 2460 8100 3420 8460
rect -5238 -780 -2276 -82
rect -5238 -1100 -5204 -780
rect -4884 -840 -2276 -780
rect -4884 -1040 -2514 -840
rect -2314 -1040 -2276 -840
rect -4884 -1100 -2276 -1040
rect -5238 -1408 -2276 -1100
rect 5344 -185 8884 -100
rect 5344 -316 8893 -185
rect 5344 -600 8168 -316
rect 5344 -1050 5550 -600
rect 6000 -950 8168 -600
rect 8820 -950 8893 -316
rect 6000 -1050 8893 -950
rect 5344 -1061 8893 -1050
rect 5344 -1370 8884 -1061
rect -1320 -9120 -360 -8760
rect -1320 -9900 -1140 -9120
rect -480 -9900 -360 -9120
rect -1320 -12840 -360 -9900
rect -1320 -13320 -1200 -12840
rect -480 -13320 -360 -12840
rect -1320 -13560 -360 -13320
rect 2400 -9120 3360 -8760
rect 2400 -9900 2580 -9120
rect 3240 -9900 3360 -9120
rect 2400 -12840 3360 -9900
rect 2400 -13320 2520 -12840
rect 3240 -13320 3360 -12840
rect 2400 -13560 3360 -13320
<< via4 >>
rect -1140 12180 -420 12660
rect 2580 12180 3300 12660
rect -5204 -1100 -4884 -780
rect 8168 -950 8820 -316
rect -1200 -13320 -480 -12840
rect 2520 -13320 3240 -12840
<< metal5 >>
rect -28066 20160 -12066 25780
rect -28066 18900 -300 20160
rect 15120 20100 31120 25800
rect 14160 20084 31120 20100
rect 2392 18968 31120 20084
rect 2392 18952 5438 18968
rect 14160 18960 31120 18968
rect -28066 17000 -12066 18900
rect -28200 16000 -12060 17000
rect -28066 9580 -12066 16000
rect -1274 13080 -306 18900
rect -1294 12660 -284 13080
rect -1294 12180 -1140 12660
rect -420 12180 -284 12660
rect -1294 11980 -284 12180
rect 2426 12660 3436 18952
rect 2426 12180 2580 12660
rect 3300 12180 3436 12660
rect 2426 11980 3436 12180
rect 15120 9600 31120 18960
rect -28000 -86 -12000 7100
rect 15030 54 31030 7066
rect -28000 -90 -4910 -86
rect -28000 -780 -4852 -90
rect -28000 -1100 -5204 -780
rect -4884 -1100 -4852 -780
rect -28000 -1376 -4852 -1100
rect 8000 -316 31030 54
rect 8000 -950 8168 -316
rect 8820 -950 31030 -316
rect -28000 -9100 -12000 -1376
rect 8000 -1486 31030 -950
rect 15030 -9134 31030 -1486
rect -28080 -19776 -12080 -11622
rect -1354 -12840 -344 -12640
rect -1354 -13320 -1200 -12840
rect -480 -13320 -344 -12840
rect -1354 -13740 -344 -13320
rect 2366 -12840 3376 -12640
rect 2366 -13320 2520 -12840
rect 3240 -13320 3376 -12840
rect -1334 -19776 -366 -13740
rect 2366 -19612 3376 -13320
rect 2332 -19628 5378 -19612
rect 15030 -19628 31030 -11764
rect -28080 -20702 -326 -19776
rect -28080 -27822 -12080 -20702
rect 2332 -20744 31030 -19628
rect 15002 -20852 31030 -20744
rect 15030 -27964 31030 -20852
<< glass >>
rect -27600 9800 -12466 25380
rect 15520 10000 30600 25400
rect -27600 -8700 -12400 6700
rect 15430 -8734 30630 6666
rect -27680 -27400 -12480 -12020
rect 15430 -27564 30630 -12164
<< end >>
