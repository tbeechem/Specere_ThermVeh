* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

sky130_fd_pr__nfet_g5v0d10v5_R72FWE a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt GSense_nFET_10VD_5Vg_1nf VD_H  VLow_Src VSUBS
XXM1 VLow_Src VSUBS VD_H sky130_fd_pr__nfet_g5v0d10v5_R72FWE
.ends

.subckt GSense_Contacts_nFT_g5_10Vd_1nf VSUBS
XGSense_nFET_10VD_5Vg_1nf_0 GSense_nFET_10VD_5Vg_1nf_0/VD_H 
+ GSense_nFET_10VD_5Vg_1nf_0/VLow_Src VSUBS GSense_nFET_10VD_5Vg_1nf
.ends

sky130_fd_pr__nfet_01v8_J36GRF a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt GSense_nFET_1f1WL150n_V1 VD_H VG_H VLow_Src 
XXM3 VD_H VG_H VLow_Src sky130_fd_pr__nfet_01v8_J36GRF
.ends

.subckt GSense_nFET_1W015L_1F_Contacts GSense_nFET_1f1WL150n_V1_0/VG_H 
XGSense_nFET_1f1WL150n_V1_0 GSense_nFET_1f1WL150n_V1_0/VD_H GSense_nFET_1f1WL150n_V1_0/VG_H
+ GSense_nFET_1f1WL150n_V1_0/VLow_Src  GSense_nFET_1f1WL150n_V1
.ends

sky130_fd_pr__nfet_03v3_nvt_XW2EXC a_n4524_n42# a_3638_n42# a_n3538_n42# a_n1764_n42#
+ a_5746_n130# a_n3914_n130# a_n3638_n130# a_6240_n42# a_n778_n42# a_2100_n42# a_50_n42#
+ a_3480_n42# a_n6950_n130# a_878_n42# a_n6674_n130# a_n5352_n42# a_n6398_n130# a_n4366_n42#
+ a_n1212_n42# a_4466_n42# a_n1982_n130# a_n2592_n42# a_3814_n130# a_3538_n130# a_n4800_n42#
+ a_n226_n42# a_n3814_n42# a_3914_n42# a_n1706_n130# a_326_n42# a_6850_n130# a_2928_n42#
+ a_n6180_n42# a_6574_n130# a_n4742_n130# a_n5194_n42# a_n2040_n42# a_5294_n42# a_6298_n130#
+ a_1882_n130# a_1154_n42# a_n1054_n42# a_n4466_n130# a_6516_n42# a_n4642_n42# a_4742_n42#
+ a_1606_n130# a_1982_n42# a_3756_n42# a_n1882_n42# a_168_n42# a_502_n130# a_n5628_n42#
+ a_4642_n130# a_n2868_n42# a_n502_n42# a_226_n130# a_602_n42# a_4366_n130# a_n2810_n130#
+ a_n2534_n130# a_996_n42# a_5570_n42# a_n2258_n130# a_n5470_n42# a_3204_n42# a_n1330_n42#
+ a_1430_n42# a_4584_n42# a_n602_n130# a_n5570_n130# a_n326_n130# a_n6456_n42# a_n5294_n130#
+ a_n3696_n42# a_n2316_n42# a_2710_n130# a_444_n42# a_2434_n130# a_n5904_n42# a_n5018_n130#
+ a_2158_n130# a_n4918_n42# a_4032_n42# a_5470_n130# a_1272_n42# a_5018_n42# a_5194_n130#
+ a_n3144_n42# a_6398_n42# a_n6298_n42# a_2258_n42# a_n3362_n130# a_n2158_n42# a_4860_n42#
+ a_n3086_n130# a_n6732_n42# a_n5746_n42# a_n384_n42# a_5846_n42# a_n3972_n42# a_n1606_n42#
+ a_1706_n42# a_n2986_n42# a_720_n42# a_n6122_n130# a_3086_n42# a_3262_n130# a_n1430_n130#
+ a_n1154_n130# a_n3420_n42# a_6674_n42# a_n6574_n42# a_4308_n42# a_n2434_n42# a_2534_n42#
+ a_5688_n42# a_1548_n42# a_n4190_n130# a_n660_n42# a_6022_n130# a_1330_n130# a_6122_n42#
+ a_1054_n130# a_778_n130# a_n6022_n42# a_5136_n42# a_n3262_n42# a_3362_n42# a_2376_n42#
+ a_n7008_n42# a_4090_n130# a_4918_n130# a_n4248_n42# a_6950_n42# a_n6850_n42# a_n2710_n42#
+ a_n1488_n42# a_2810_n42# a_5964_n42# a_n878_n130# a_1824_n42# a_n108_n42# a_n4090_n42#
+ a_4190_n42# a_n5846_n130# a_2986_n130# a_n50_n130# a_n5076_n42# a_n936_n42# a_5412_n42#
+ a_6792_n42# a_2652_n42# a_n7142_n264# m1_n6988_n248#
X0 a_n6022_n42# a_n6122_n130# a_n6180_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1 a_n3538_n42# a_n3638_n130# a_n3696_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X2 a_3086_n42# a_2986_n130# a_2928_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X3 a_6950_n42# a_6850_n130# a_6792_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X4 a_n3262_n42# a_n3362_n130# a_n3420_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X5 a_5294_n42# a_5194_n130# a_5136_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X6 a_6674_n42# a_6574_n130# a_6516_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X7 a_n4642_n42# a_n4742_n130# a_n4800_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X8 a_n2986_n42# a_n3086_n130# a_n3144_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X9 a_1706_n42# a_1606_n130# a_1548_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X10 a_6398_n42# a_6298_n130# a_6240_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X11 a_n4366_n42# a_n4466_n130# a_n4524_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X12 a_n1882_n42# a_n1982_n130# a_n2040_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X13 a_n502_n42# a_n602_n130# a_n660_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X14 a_1430_n42# a_1330_n130# a_1272_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X15 a_50_n42# a_n50_n130# a_n108_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X16 a_n5746_n42# a_n5846_n130# a_n5904_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X17 a_2810_n42# a_2710_n130# a_2652_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X18 a_n4090_n42# a_n4190_n130# a_n4248_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X19 a_878_n42# a_778_n130# a_720_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X20 a_1154_n42# a_1054_n130# a_996_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X21 a_n226_n42# a_n326_n130# a_n384_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X22 a_n5470_n42# a_n5570_n130# a_n5628_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X23 a_2534_n42# a_2434_n130# a_2376_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X24 a_n5194_n42# a_n5294_n130# a_n5352_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X25 a_n6850_n42# a_n6950_n130# a_n7008_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X26 a_2258_n42# a_2158_n130# a_2100_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X27 a_3914_n42# a_3814_n130# a_3756_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X28 a_6122_n42# a_6022_n130# a_5964_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X29 a_n6574_n42# a_n6674_n130# a_n6732_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X30 a_3638_n42# a_3538_n130# a_3480_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X31 a_n1606_n42# a_n1706_n130# a_n1764_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X32 a_n6298_n42# a_n6398_n130# a_n6456_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X33 a_3362_n42# a_3262_n130# a_3204_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X34 a_5018_n42# a_4918_n130# a_4860_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X35 a_602_n42# a_502_n130# a_444_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X36 a_n1330_n42# a_n1430_n130# a_n1488_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X37 a_4742_n42# a_4642_n130# a_4584_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X38 a_n2710_n42# a_n2810_n130# a_n2868_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X39 a_n1054_n42# a_n1154_n130# a_n1212_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X40 a_326_n42# a_226_n130# a_168_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X41 a_1982_n42# a_1882_n130# a_1824_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X42 a_4466_n42# a_4366_n130# a_4308_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X43 a_n4918_n42# a_n5018_n130# a_n5076_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X44 a_n2434_n42# a_n2534_n130# a_n2592_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X45 a_4190_n42# a_4090_n130# a_4032_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X46 a_5846_n42# a_5746_n130# a_5688_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X47 a_n3814_n42# a_n3914_n130# a_n3972_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X48 a_n2158_n42# a_n2258_n130# a_n2316_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X49 a_n778_n42# a_n878_n130# a_n936_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X50 a_5570_n42# a_5470_n130# a_5412_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
.ends

sky130_fd_pr__nfet_03v3_nvt_XW2EXC
.subckt GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH VG_H  VLow_Src li_174_n490# VSUBS
XXM1 VLow_Src VD_H VLow_Src VLow_Src VG_H VG_H VG_H VLow_Src VD_H VD_H VLow_Src VLow_Src
+ li_174_n490# VD_H VG_H VD_H VG_H VD_H VLow_Src VLow_Src VG_H VD_H VG_H VG_H VD_H
+ VD_H VD_H VLow_Src VG_H VD_H VG_H VLow_Src VLow_Src VG_H VG_H VLow_Src VD_H VD_H
+ VG_H VG_H VLow_Src VD_H VG_H VD_H VLow_Src VD_H VG_H VD_H VD_H VLow_Src VLow_Src
+ VG_H VLow_Src VG_H VLow_Src VLow_Src VG_H VLow_Src VG_H VG_H VG_H VD_H VLow_Src
+ VG_H VD_H VD_H VLow_Src VD_H VLow_Src VG_H VG_H VG_H VD_H VG_H VD_H VLow_Src VG_H
+ VD_H VG_H VD_H VG_H VG_H VD_H VLow_Src VG_H VLow_Src VLow_Src VG_H VD_H VD_H VLow_Src
+ VLow_Src VG_H VD_H VD_H VG_H VLow_Src VLow_Src VLow_Src VD_H VLow_Src VD_H VLow_Src
+ VLow_Src VLow_Src VG_H VD_H VG_H VG_H VG_H VLow_Src VLow_Src VD_H VD_H VLow_Src
+ VD_H VLow_Src VD_H VG_H VD_H VG_H VG_H VLow_Src VG_H VG_H VD_H VLow_Src VD_H VLow_Src
+ VLow_Src VD_H VG_H VG_H VD_H VD_H VLow_Src VD_H VD_H VLow_Src VD_H VG_H VLow_Src
+ VD_H VLow_Src VD_H VG_H VG_H VG_H VLow_Src VLow_Src VD_H VLow_Src VD_H VSUBS VD_H
.ends

.subckt nFET_3p3Vd_3VG_51NF_LTherm_Contacts  VSUBS
XGSense_nFET_3VD_3Vg_51nf_V2AllGates_VH_0 GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH_0/VG_H
+  GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH_0/VLow_Src
+ m1_n4654_560# VSUBS GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH
.ends

sky130_fd_pr__nfet_03v3_nvt_XW2EXC
.subckt GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline VG_H  VLow_Src m1_6800_n480#
+ VSUBS
XXM1 VLow_Src VD_H VLow_Src VLow_Src VG_H VG_H VG_H VLow_Src VD_H VD_H VLow_Src VLow_Src
+ VG_H VD_H VG_H VD_H VG_H VD_H VLow_Src VLow_Src VG_H VD_H VG_H VG_H VD_H VD_H VD_H
+ VLow_Src VG_H VD_H VG_H VLow_Src VLow_Src VG_H VG_H VLow_Src VD_H VD_H VG_H VG_H
+ VLow_Src VD_H VG_H VD_H VLow_Src VD_H VG_H VD_H VD_H VLow_Src VLow_Src VG_H VLow_Src
+ VG_H VLow_Src VLow_Src VG_H VLow_Src VG_H VG_H VG_H VD_H VLow_Src VG_H VD_H VD_H
+ VLow_Src VD_H VLow_Src VG_H VG_H m1_6800_n480# VD_H VG_H VD_H VLow_Src VG_H VD_H
+ VG_H VD_H VG_H VG_H VD_H VLow_Src VG_H VLow_Src VLow_Src VG_H VD_H VD_H VLow_Src
+ VLow_Src VG_H VD_H VD_H VG_H VLow_Src VLow_Src VLow_Src VD_H VLow_Src VD_H VLow_Src
+ VLow_Src VLow_Src VG_H VD_H VG_H VG_H VG_H VLow_Src VLow_Src VD_H VD_H VLow_Src
+ VD_H VLow_Src VD_H VG_H VD_H VG_H VG_H VLow_Src VG_H VG_H VD_H VLow_Src VD_H VLow_Src
+ VLow_Src VD_H VG_H VG_H VD_H VD_H VLow_Src VD_H VD_H VLow_Src VD_H VG_H VLow_Src
+ VD_H VLow_Src VD_H VG_H VG_H VG_H VLow_Src VLow_Src VD_H VLow_Src VD_H VSUBS VD_H
.ends

.subckt nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts  VSUBS
XGSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0 GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0/VG_H
+  GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline_0/VLow_Src
+ m2_n1290_6370# VSUBS GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_W5U4AW c2_n3079_n3000# m4_n3179_n3100#
X0 c2_n3079_n3000# m4_n3179_n3100# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
.ends

.subckt sky130_fd_sc_hvl__buf_8 VPWR   VGND X A
X0 X a_45_443# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5 M=8
X1 X a_45_443# VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5 M=8
X2 a_45_443# A VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.2025 ps=1.29 w=0.75 l=0.5 M=3
X3 VPWR A a_45_443# sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5 M=3
.ends

sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ a_n683_n200# a_n189_n297# a_29_n297# a_189_n200#
+ a_n901_n200# a_247_n297# a_n407_n297# a_465_n297# a_407_n200# a_n625_n297# a_683_n297#
+ a_625_n200# a_n843_n297# w_n1101_n497# a_843_n200# a_n29_n200# a_n247_n200# a_n465_n200#
X0 a_n247_n200# a_n407_n297# a_n465_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X1 a_843_n200# a_683_n297# a_625_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X2 a_407_n200# a_247_n297# a_189_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X3 a_189_n200# a_29_n297# a_n29_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X4 a_n465_n200# a_n625_n297# a_n683_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X5 a_625_n200# a_465_n297# a_407_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X6 a_n29_n200# a_n189_n297# a_n247_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X7 a_n683_n200# a_n843_n297# a_n901_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
.ends

sky130_fd_pr__nfet_g5v0d10v5_TGFUGS a_n792_n200# a_298_n200# a_516_n200# a_734_n200#
+ a_n926_n422# a_138_n288# a_n298_n288# a_80_n200# a_356_n288# a_n516_n288# a_574_n288#
+ a_n734_n288# a_n138_n200# a_n356_n200# a_n574_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X1 a_n574_n200# a_n734_n288# a_n792_n200# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
X2 a_734_n200# a_574_n288# a_516_n200# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X3 a_298_n200# a_138_n288# a_80_n200# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X4 a_n138_n200# a_n298_n288# a_n356_n200# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X5 a_n356_n200# a_n516_n288# a_n574_n200# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X6 a_516_n200# a_356_n288# a_298_n200# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
.ends

sky130_fd_pr__res_xhigh_po_0p69_S5N9F3 a_124_2496# a_n4122_n2932# a_n4122_2496#
+ a_2054_n2932# a_2054_2496# a_896_n2932# a_510_2496# a_3598_2496# a_3984_2496# a_3598_n2932#
+ a_2440_2496# a_n3736_n2932# a_1668_n2932# a_n1806_n2932# a_5142_n2932# a_510_n2932#
+ a_n2192_2496# a_n3736_2496# a_3212_n2932# a_n5410_n3062# a_1668_2496# a_n262_2496#
+ a_4756_n2932# a_5142_2496# a_2826_n2932# a_n2192_n2932# a_n1806_2496# a_n5280_2496#
+ a_n648_n2932# a_n5280_n2932# a_n3350_n2932# a_4756_2496# a_3212_2496# a_1282_n2932#
+ a_124_n2932# a_n1420_n2932# a_n4894_n2932# a_896_2496# a_n2964_n2932# a_n3350_2496#
+ a_n4508_2496# a_n4894_2496# a_n4508_n2932# a_4370_n2932# a_1282_2496# a_2826_2496#
+ a_2440_n2932# a_3984_n2932# a_n1034_2496# a_n2578_2496# a_n1420_2496# a_n2964_2496#
+ a_n262_n2932# a_n648_2496# a_n1034_n2932# a_4370_2496# a_n2578_n2932#
X0 a_n262_2496# a_n262_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X1 a_n3350_2496# a_n3350_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X2 a_n4122_2496# a_n4122_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X3 a_n4894_2496# a_n4894_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X4 a_n3736_2496# a_n3736_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X5 a_1282_2496# a_1282_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X6 a_5142_2496# a_5142_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X7 a_4756_2496# a_4756_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X8 a_124_2496# a_124_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X9 a_510_2496# a_510_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X10 a_896_2496# a_896_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X11 a_n5280_2496# a_n5280_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X12 a_n648_2496# a_n648_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X13 a_n4508_2496# a_n4508_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X14 a_n2192_2496# a_n2192_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X15 a_n1034_2496# a_n1034_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X16 a_2054_2496# a_2054_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X17 a_1668_2496# a_1668_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X18 a_2440_2496# a_2440_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X19 a_n1420_2496# a_n1420_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X20 a_n2578_2496# a_n2578_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X21 a_n1806_2496# a_n1806_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X22 a_3212_2496# a_3212_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X23 a_3598_2496# a_3598_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X24 a_n2964_2496# a_n2964_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X25 a_4370_2496# a_4370_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X26 a_2826_2496# a_2826_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
X27 a_3984_2496# a_3984_n2932# sky130_fd_pr__res_xhigh_po_0p69 l=25.12
.ends

sky130_fd_pr__pfet_g5v0d10v5_3YBPVB a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_sc_hvl__schmittbuf_1 X A   VPWR VGND
X0 X a_117_181# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.315925 ps=1.45 w=0.75 l=0.5
X1 a_217_207# a_117_181# a_64_207# sky130_fd_pr__nfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.5
X2 VPWR A a_231_463# sky130_fd_pr__pfet_g5v0d10v5 ad=0.34075 pd=1.73 as=0.105 ps=1.03 w=0.75 l=0.5
X3 VGND A a_217_207# sky130_fd_pr__nfet_g5v0d10v5 ad=0.315925 pd=1.45 as=0.0588 ps=0.7 w=0.42 l=0.5
X4 a_78_463# VGND sky130_fd_pr__res_generic_nd__hv w=0.29 l=1.355
X5 a_64_207# VPWR sky130_fd_pr__res_generic_pd__hv w=0.29 l=3.11
X6 X a_117_181# VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.34075 ps=1.73 w=1.5 l=0.5
X7 a_231_463# A a_117_181# sky130_fd_pr__pfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X8 a_231_463# a_117_181# a_78_463# sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X9 a_217_207# A a_117_181# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.5
.ends

sky130_fd_pr__pfet_g5v0d10v5_YUHPXE a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

sky130_fd_pr__nfet_g5v0d10v5_PKVMTM a_80_n200# a_n272_n422# a_n138_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC a_80_n200# a_n272_n422# a_n138_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_WRT4AW c1_n3036_n3000# m3_n3136_n3100#
X0 c1_n3036_n3000# m3_n3136_n3100# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
.ends

sky130_fd_pr__pfet_g5v0d10v5_YEUEBV a_n792_n200# a_138_n297# a_n298_n297#
+ a_298_n200# a_356_n297# a_n516_n297# a_574_n297# a_516_n200# a_n734_n297# a_734_n200#
+ a_n80_n297# a_80_n200# a_n138_n200# a_n356_n200# a_n574_n200# w_n992_n497#
X0 a_80_n200# a_n80_n297# a_n138_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X1 a_n574_n200# a_n734_n297# a_n792_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
X2 a_734_n200# a_574_n297# a_516_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X3 a_298_n200# a_138_n297# a_80_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X4 a_n138_n200# a_n298_n297# a_n356_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X5 a_n356_n200# a_n516_n297# a_n574_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X6 a_516_n200# a_356_n297# a_298_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
.ends

sky130_fd_pr__pfet_g5v0d10v5_YUHPBG a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_sc_hvl__inv_8  VGND VPWR  Y A
X0 Y A VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5 M=8
X1 VGND A Y sky130_fd_pr__nfet_g5v0d10v5 ad=0.1575 pd=1.17 as=0.105 ps=1.03 w=0.75 l=0.5 M=8
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__fill_4 abstract view
.subckt sky130_fd_sc_hvl__fill_4    
.ends

sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
.subckt example_por vdd3v3 vdd1v8 vss porb_h por_l porb_l
Xsky130_fd_pr__cap_mim_m3_2_W5U4AW_0 vss sky130_fd_sc_hvl__schmittbuf_1_0/A sky130_fd_pr__cap_mim_m3_2_W5U4AW
Xsky130_fd_sc_hvl__buf_8_1 vdd1v8   vss porb_l sky130_fd_sc_hvl__inv_8_0/A
+ sky130_fd_sc_hvl__buf_8
Xsky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ_0 m1_502_7653# m1_502_7653# m1_502_7653# m1_502_7653#
+ vdd3v3 m1_502_7653# m1_502_7653# m1_502_7653# vdd3v3 m1_502_7653# m1_502_7653# m1_502_7653#
+ m1_502_7653# vdd3v3 vdd3v3 vdd3v3 m1_502_7653# sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ
Xsky130_fd_pr__nfet_g5v0d10v5_TGFUGS_0 m1_721_6815# vss m1_721_6815# vss vss m1_721_6815#
+ m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# vss
+ m1_721_6815# vss sky130_fd_pr__nfet_g5v0d10v5_TGFUGS
Xsky130_fd_pr__res_xhigh_po_0p69_S5N9F3_0 li_5638_5813# li_1391_165# li_1006_5813#
+ li_7567_165# li_7182_5813# li_6023_165# li_5638_5813# li_8726_5813# li_9498_5813#
+ li_9111_165# li_7954_5813# li_1391_165# li_6795_165# li_3707_165# vss li_6023_165#
+ li_3322_5813# li_1778_5813# li_8339_165# vss li_7182_5813# li_4866_5813# li_9883_165#
+ vss li_8339_165# li_2935_165# li_3322_5813# vss li_4479_165# vss li_2163_165# vdd3v3
+ li_8726_5813# li_6795_165# li_5251_165# li_3707_165# li_619_165# li_6410_5813# li_2163_165#
+ li_1778_5813# li_1006_5813# vss li_619_165# li_9883_165# li_6410_5813# li_7954_5813#
+ li_7567_165# li_9111_165# li_4094_5813# li_2550_5813# li_4094_5813# li_2550_5813#
+ li_5251_165# li_4866_5813# li_4479_165# li_9498_5813# sky130_fd_pr__res_xhigh_po_0p69_S5N9F3
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_0 m1_2756_6573# sky130_fd_sc_hvl__schmittbuf_1_0/A
+ vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_sc_hvl__schmittbuf_1_0 sky130_fd_sc_hvl__inv_8_0/A sky130_fd_sc_hvl__schmittbuf_1_0/A
+   vdd3v3 vss sky130_fd_sc_hvl__schmittbuf_1
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_1 m1_185_6573# m1_721_6815# vdd3v3 m1_2993_7658#
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_2 m1_2756_6573# m1_4283_8081# vdd3v3 m1_2756_6573#
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_3 m1_185_6573# m1_502_7653# vdd3v3 m1_185_6573#
Xsky130_fd_pr__pfet_g5v0d10v5_YUHPXE_0 m1_4283_8081# m1_6249_7690# vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_YUHPXE
Xsky130_fd_pr__nfet_g5v0d10v5_PKVMTM_0 m1_2756_6573# vss vss sky130_fd_pr__nfet_g5v0d10v5_PKVMTM
Xsky130_fd_pr__nfet_g5v0d10v5_ZK8HQC_0 m1_185_6573# vss vss sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC
Xsky130_fd_pr__cap_mim_m3_1_WRT4AW_0 sky130_fd_sc_hvl__schmittbuf_1_0/A vss sky130_fd_pr__cap_mim_m3_1_WRT4AW
Xsky130_fd_pr__pfet_g5v0d10v5_YEUEBV_0 vdd3v3 m1_4283_8081# m1_4283_8081# m1_4283_8081#
+ m1_4283_8081# m1_4283_8081# m1_4283_8081# vdd3v3 m1_4283_8081# m1_4283_8081# m1_4283_8081#
+ vdd3v3 m1_4283_8081# vdd3v3 m1_4283_8081# sky130_fd_pr__pfet_g5v0d10v5_YEUEBV
Xsky130_fd_pr__pfet_g5v0d10v5_YUHPBG_0 m1_502_7653# m1_2993_7658# vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_YUHPBG
Xsky130_fd_sc_hvl__inv_8_0  vss vdd1v8  por_l sky130_fd_sc_hvl__inv_8_0/A
+ sky130_fd_sc_hvl__inv_8
Xsky130_fd_sc_hvl__buf_8_0 vdd3v3   vss porb_h sky130_fd_sc_hvl__inv_8_0/A
+ sky130_fd_sc_hvl__buf_8
.ends

.subckt user_analog_proj_example example_por_0/por_l example_por_1/por_l example_por_0/vdd1v8
+ example_por_1/vdd3v3 example_por_1/porb_l example_por_0/vdd3v3 example_por_1/porb_h
+ example_por_0/porb_l example_por_0/porb_h VSUBS example_por_1/vdd1v8
Xexample_por_0 example_por_0/vdd3v3 example_por_0/vdd1v8 VSUBS example_por_0/porb_h
+ example_por_0/por_l example_por_0/porb_l example_por
Xexample_por_1 example_por_1/vdd3v3 example_por_1/vdd1v8 VSUBS example_por_1/porb_h
+ example_por_1/por_l example_por_1/porb_l example_por
.ends

sky130_fd_pr__pfet_g5v0d10v5_WLCVX2 a_n50_n197# a_50_n100# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt GSense_pFET_10VD_5Vg_1nf  VLow_Src VG_H
XXM1 VG_H VLow_Src sky130_fd_pr__pfet_g5v0d10v5_WLCVX2
.ends

.subckt GSense_pFET_10Vd_5p5Vg_1nf
XGSense_pFET_10VD_5Vg_1nf_0  GSense_pFET_10VD_5Vg_1nf_0/VLow_Src
+ GSense_pFET_10VD_5Vg_1nf_0/VG_H GSense_pFET_10VD_5Vg_1nf
.ends

sky130_fd_pr__nfet_03v3_nvt_J2JJF2 a_858_n42# a_30_n42# a_306_n42# a_n798_n42#
+ a_n1292_n130# a_1134_n42# a_n1016_n130# a_n246_n42# a_1192_n130# a_n1074_n42# a_916_n130#
+ a_n1484_n264# a_188_n42# a_n522_n42# a_n1350_n42# a_n88_n42# a_464_n42# a_n364_n42#
+ a_1292_n42# a_n1192_n42# a_n640_n42# a_740_n42# a_582_n42# a_640_n130# a_364_n130#
+ a_88_n130# a_n740_n130# a_1016_n42# a_n916_n42# a_n188_n130# a_n464_n130#
X0 a_740_n42# a_640_n130# a_582_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1 a_n1192_n42# a_n1292_n130# a_n1350_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X2 a_464_n42# a_364_n130# a_306_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X3 a_n916_n42# a_n1016_n130# a_n1074_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X4 a_188_n42# a_88_n130# a_30_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X5 a_n640_n42# a_n740_n130# a_n798_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X6 a_1292_n42# a_1192_n130# a_1134_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X7 a_n364_n42# a_n464_n130# a_n522_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X8 a_n88_n42# a_n188_n130# a_n246_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X9 a_1016_n42# a_916_n130# a_858_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
.ends

.subckt GSense_nFET_3VD_3Vg_10nf_V2 VG_H VD_H VLow_Src m1_1152_n620# VSUBS
XXM1 VD_H VLow_Src VD_H VD_H VG_H VLow_Src VG_H VD_H VG_H VLow_Src VG_H VSUBS VD_H
+ VLow_Src VD_H VLow_Src VLow_Src VD_H VD_H VLow_Src VLow_Src VD_H VLow_Src VG_H VG_H
+ VG_H VG_H VLow_Src VD_H m1_1152_n620# sky130_fd_pr__nfet_03v3_nvt_J2JJF2
.ends

.subckt nFET_3VD_3VG_10nF_Contacts  VSUBS
XGSense_nFET_3VD_3Vg_10nf_V2_0 GSense_nFET_3VD_3Vg_10nf_V2_0/VG_H GSense_nFET_3VD_3Vg_10nf_V2_0/VD_H
+ GSense_nFET_3VD_3Vg_10nf_V2_0/VLow_Src m1_n1260_1140# VSUBS GSense_nFET_3VD_3Vg_10nf_V2
.ends

sky130_fd_pr__nfet_03v3_nvt_EJ4KLV a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# sky130_fd_pr__nfet_03v3_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt GSense_nFET_3VD_3Vg_1nf VD_H  VLow_Src VSUBS
XXM1 VLow_Src VSUBS VD_H sky130_fd_pr__nfet_03v3_nvt_EJ4KLV
.ends

.subckt GSense_Contacts_nFET_3V_1nf VSUBS
XGSense_nFET_3VD_3Vg_1nf_0 GSense_nFET_3VD_3Vg_1nf_0/VD_H 
+ GSense_nFET_3VD_3Vg_1nf_0/VLow_Src VSUBS GSense_nFET_3VD_3Vg_1nf
.ends

.subckt nFET_3VD_3VG_50nF_Therm_FET12  VSUBS
XGSense_nFET_3VD_3Vg_51nf_V2AllGates_Mid_Therm_0 GSense_nFET_3VD_3Vg_51nf_V2AllGates_Mid_Therm_0/VG_H
+  GSense_nFET_3VD_3Vg_51nf_V2AllGates_Mid_Therm_0/VLow_Src
+ m2_n1312_3142# VSUBS GSense_nFET_3VD_3Vg_51nf_V2AllGates_Therm_Midline
.ends

sky130_fd_pr__nfet_03v3_nvt_VB5P9F a_50_n42# a_326_n42# a_n226_n42# a_168_n42#
+ a_502_n130# a_602_n42# a_n502_n42# a_226_n130# a_n602_n130# a_n326_n130# a_444_n42#
+ a_n794_n264# a_n384_n42# a_n660_n42# a_n108_n42# a_n50_n130#
X0 a_n502_n42# a_n602_n130# a_n660_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1 a_50_n42# a_n50_n130# a_n108_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X2 a_n226_n42# a_n326_n130# a_n384_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X3 a_602_n42# a_502_n130# a_444_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X4 a_326_n42# a_226_n130# a_168_n42# sky130_fd_pr__nfet_03v3_nvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
.ends

.subckt GSense_nFET_3VD_3Vg_5nf_V2 VD_H VG_H VLow_Src  VSUBS
Xsky130_fd_pr__nfet_03v3_nvt_VB5P9F_0 VLow_Src VD_H VD_H VLow_Src VG_H VLow_Src VLow_Src
+ VG_H VG_H VG_H VD_H VSUBS VLow_Src VD_H VD_H sky130_fd_pr__nfet_03v3_nvt_VB5P9F
.ends

.subckt GSense_nFET_3p3V_5nF_Contacts_V2 VSUBS
XGSense_nFET_3VD_3Vg_5nf_V2_1 GSense_nFET_3VD_3Vg_5nf_V2_1/VD_H GSense_nFET_3VD_3Vg_5nf_V2_1/VG_H
+ GSense_nFET_3VD_3Vg_5nf_V2_1/VLow_Src  VSUBS GSense_nFET_3VD_3Vg_5nf_V2
.ends

sky130_fd_pr__pfet_01v8_8JS3FC a_n73_n100# a_15_n100# a_n33_n197#
X0 a_15_n100# a_n33_n197# a_n73_n100# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt GSense_pFET_1p8VD_1p8Vg_1nf VD_H VLow_Src 
XXM1 VD_H VLow_Src sky130_fd_pr__pfet_01v8_8JS3FC
.ends

.subckt GSense_Contacts_pfet_1p8Vd_1p8Vg
XGSense_pFET_1p8VD_1p8Vg_1nf_0 GSense_pFET_1p8VD_1p8Vg_1nf_0/VD_H GSense_pFET_1p8VD_1p8Vg_1nf_0/VLow_Src
+  GSense_pFET_1p8VD_1p8Vg_1nf
.ends

.subckt user_project_wrapper    
+   gpio_analog[3]   
+ gpio_analog[7]     
+  io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2]     
+ io_oeb[11] io_oeb[12]   io_oeb[15] io_oeb[16]  
+    io_out[11] io_out[12]   io_out[15]
+ io_out[16]       
+ vccd1          
+      io_analog[4]_uq3
+  vssa1_uq1      
+ vdda1_uq1 vssd1
XGSense_Contacts_nFT_g5_10Vd_1nf_1 vssa1_uq1 GSense_Contacts_nFT_g5_10Vd_1nf
XGSense_Contacts_nFT_g5_10Vd_1nf_2 vssa1_uq1 GSense_Contacts_nFT_g5_10Vd_1nf
XGSense_nFET_1W015L_1F_Contacts_0 GSense_nFET_1W015L_1F_Contacts_0/GSense_nFET_1f1WL150n_V1_0/VG_H
+  GSense_nFET_1W015L_1F_Contacts
XGSense_nFET_1W015L_1F_Contacts_2 GSense_nFET_1W015L_1F_Contacts_2/GSense_nFET_1f1WL150n_V1_0/VG_H
+  GSense_nFET_1W015L_1F_Contacts
XGSense_nFET_1W015L_1F_Contacts_1 GSense_nFET_1W015L_1F_Contacts_1/GSense_nFET_1f1WL150n_V1_0/VG_H
+  GSense_nFET_1W015L_1F_Contacts
XGSense_nFET_1W015L_1F_Contacts_3 GSense_nFET_1W015L_1F_Contacts_3/GSense_nFET_1f1WL150n_V1_0/VG_H
+  GSense_nFET_1W015L_1F_Contacts
XnFET_3p3Vd_3VG_51NF_LTherm_Contacts_0 
+ vssa1_uq1 nFET_3p3Vd_3VG_51NF_LTherm_Contacts
XnFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_0 
+ vssa1_uq1 nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts
XnFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_1 
+ vssa1_uq1 nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts
XnFET_3p3Vd_3VG_51NF_LTherm_Contacts_1  vssa1_uq1 nFET_3p3Vd_3VG_51NF_LTherm_Contacts
XGSense_nFET_1W015L_1F_Contacts_4 GSense_nFET_1W015L_1F_Contacts_4/GSense_nFET_1f1WL150n_V1_0/VG_H
+  GSense_nFET_1W015L_1F_Contacts
Xuser_analog_proj_example_0 io_out[16] io_out[12] vccd1 vdda1_uq1 io_out[11] io_analog[4]_uq3
+ gpio_analog[3] io_out[15] gpio_analog[7] vssa1_uq1 vccd1 user_analog_proj_example
XnFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_2 
+ vssa1_uq1 nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts
XnFET_3p3Vd_3VG_51NF_LTherm_Contacts_2 
+ vssa1_uq1 nFET_3p3Vd_3VG_51NF_LTherm_Contacts
XGSense_nFET_1W015L_1F_Contacts_5 GSense_nFET_1W015L_1F_Contacts_5/GSense_nFET_1f1WL150n_V1_0/VG_H
+  GSense_nFET_1W015L_1F_Contacts
XnFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_3  vssa1_uq1 nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts
XnFET_3VD_3VG_50NF_MiDLine_Therm_Contacts_5 
+ vssa1_uq1 nFET_3VD_3VG_50NF_MiDLine_Therm_Contacts
XnFET_3VD_3VG_10nF_Contacts_0  vssa1_uq1
+ nFET_3VD_3VG_10nF_Contacts
XGSense_Contacts_nFET_3V_1nf_0 vssa1_uq1 GSense_Contacts_nFET_3V_1nf
XnFET_3VD_3VG_10nF_Contacts_1  vssa1_uq1
+ nFET_3VD_3VG_10nF_Contacts
XGSense_Contacts_nFET_3V_1nf_1 vssa1_uq1 GSense_Contacts_nFET_3V_1nf
XnFET_3VD_3VG_10nF_Contacts_2  vssa1_uq1
+ nFET_3VD_3VG_10nF_Contacts
XnFET_3VD_3VG_50nF_Therm_FET12_0  vssa1_uq1
+ nFET_3VD_3VG_50nF_Therm_FET12
XnFET_3VD_3VG_10nF_Contacts_3  vssa1_uq1 nFET_3VD_3VG_10nF_Contacts
XGSense_Contacts_nFET_3V_1nf_2 vssa1_uq1 GSense_Contacts_nFET_3V_1nf
XnFET_3VD_3VG_50nF_Therm_FET12_1  vssa1_uq1 nFET_3VD_3VG_50nF_Therm_FET12
XGSense_Contacts_nFET_3V_1nf_3 vssa1_uq1 GSense_Contacts_nFET_3V_1nf
XGSense_nFET_3p3V_5nF_Contacts_V2_0 vssa1_uq1 GSense_nFET_3p3V_5nF_Contacts_V2
XnFET_3VD_3VG_50nF_Therm_FET12_3  vssa1_uq1
+ nFET_3VD_3VG_50nF_Therm_FET12
XGSense_nFET_3p3V_5nF_Contacts_V2_1 vssa1_uq1 GSense_nFET_3p3V_5nF_Contacts_V2
XGSense_nFET_3p3V_5nF_Contacts_V2_2 vssa1_uq1 GSense_nFET_3p3V_5nF_Contacts_V2
XGSense_Contacts_nFT_g5_10Vd_1nf_0 vssa1_uq1 GSense_Contacts_nFT_g5_10Vd_1nf
R0 io_oeb[15] vssd1 sky130_fd_pr__res_generic_m3 w=0.56 l=0.6
R1 io_clamp_high[0] io_analog[4]_uq3 sky130_fd_pr__res_generic_m3 w=11 l=0.25
R2 vssd1 io_oeb[11] sky130_fd_pr__res_generic_m3 w=0.56 l=0.58
R3 io_clamp_low[1] vssa1_uq1 sky130_fd_pr__res_generic_m3 w=11 l=0.25
R4 io_oeb[16] vssd1 sky130_fd_pr__res_generic_m3 w=0.56 l=0.31
R5 io_clamp_low[0] vssa1_uq1 sky130_fd_pr__res_generic_m3 w=11 l=0.25
R6 vssd1 io_oeb[12] sky130_fd_pr__res_generic_m3 w=0.56 l=0.49
R7 io_clamp_high[2] vssa1_uq1 sky130_fd_pr__res_generic_m3 w=11 l=0.25
R8 io_clamp_high[1] vssa1_uq1 sky130_fd_pr__res_generic_m3 w=11 l=0.25
R9 io_clamp_low[2] vssa1_uq1 sky130_fd_pr__res_generic_m3 w=11 l=0.25
.ends

