magic
tech sky130A
magscale 1 2
timestamp 1717386517
<< metal1 >>
rect 5996 12654 7448 13018
rect 5996 11830 6392 12654
rect 7118 11830 7448 12654
rect 5996 2684 7448 11830
rect -4654 1362 -4134 1596
rect -4654 1238 -4490 1362
rect -4382 1238 -4134 1362
rect -4654 560 -4134 1238
rect -6611 -112 -6605 214
rect -6279 -112 -5742 214
rect 10392 -530 11192 394
rect 10392 -776 10462 -530
rect 10602 -776 11192 -530
rect 10392 -862 11192 -776
rect -5528 -1248 -366 -1048
rect -5528 -2650 -5204 -1248
rect -5526 -2994 -5262 -2650
rect -6088 -11910 -4636 -2994
rect -6088 -12734 -5758 -11910
rect -5032 -12734 -4636 -11910
rect -6088 -13328 -4636 -12734
<< via1 >>
rect 6392 11830 7118 12654
rect -4490 1238 -4382 1362
rect -6605 -112 -6279 214
rect -4502 -640 -4434 -584
rect 10462 -776 10602 -530
rect -5758 -12734 -5032 -11910
<< metal2 >>
rect 6030 14670 7350 15100
rect 6030 13944 6392 14670
rect 7084 13944 7350 14670
rect 6030 12654 7350 13944
rect 6030 11830 6392 12654
rect 7118 11830 7350 12654
rect 6030 11468 7350 11830
rect -1260 6240 -300 6360
rect -1260 5580 -1080 6240
rect -420 5580 -300 6240
rect -1260 4689 -300 5580
rect 2460 6240 3420 6360
rect 2460 5580 2640 6240
rect 3300 5580 3420 6240
rect 2460 4689 3420 5580
rect -3670 4674 3429 4689
rect -4664 3617 3429 4674
rect -4664 1456 -4102 3617
rect -4654 1362 -4118 1456
rect -4654 1238 -4490 1362
rect -4382 1238 -4118 1362
rect -4654 1076 -4118 1238
rect -6605 214 -6279 220
rect -7444 -112 -7435 214
rect -7109 -112 -6605 214
rect -6605 -118 -6279 -112
rect 10398 -440 11194 -438
rect 10398 -530 11393 -440
rect -4510 -584 -4428 -566
rect -4510 -640 -4502 -584
rect -4434 -640 -4428 -584
rect -4510 -1814 -4428 -640
rect 10398 -776 10462 -530
rect 10602 -776 11393 -530
rect 10398 -858 11393 -776
rect 10794 -862 11393 -858
rect 11815 -862 11824 -440
rect 2400 -1814 3360 -1812
rect -4518 -2766 3376 -1814
rect -1320 -6240 -360 -2766
rect -1320 -6900 -1140 -6240
rect -480 -6900 -360 -6240
rect -1320 -7020 -360 -6900
rect 2400 -6240 3360 -2766
rect 2400 -6900 2580 -6240
rect 3240 -6900 3360 -6240
rect 2400 -7020 3360 -6900
rect -6054 -11910 -4734 -11742
rect -6054 -12734 -5758 -11910
rect -5032 -12734 -4734 -11910
rect -6054 -14352 -4734 -12734
rect -6054 -15078 -5790 -14352
rect -5098 -15078 -4734 -14352
rect -6054 -15374 -4734 -15078
<< via2 >>
rect 6392 13944 7084 14670
rect -1080 5580 -420 6240
rect 2640 5580 3300 6240
rect -7435 -112 -7109 214
rect 11393 -862 11815 -440
rect -1140 -6900 -480 -6240
rect 2580 -6900 3240 -6240
rect -5790 -15078 -5098 -14352
<< metal3 >>
rect 6126 17284 7316 17692
rect 6126 16360 6352 17284
rect 7028 16360 7316 17284
rect 6126 14670 7316 16360
rect 6126 13944 6392 14670
rect 7084 13944 7316 14670
rect 6126 13596 7316 13944
rect -1260 9240 -300 9480
rect -1260 8460 -1080 9240
rect -420 8460 -300 9240
rect -1260 6240 -300 8460
rect -1260 5580 -1080 6240
rect -420 5580 -300 6240
rect -1260 5400 -300 5580
rect 2460 9240 3420 9480
rect 2460 8460 2640 9240
rect 3300 8460 3420 9240
rect 2460 6240 3420 8460
rect 2460 5580 2640 6240
rect 3300 5580 3420 6240
rect 2460 5400 3420 5580
rect -7440 214 -7104 219
rect -8129 -112 -8123 214
rect -7797 -112 -7435 214
rect -7109 -112 -7104 214
rect -7440 -117 -7104 -112
rect 11388 -440 11820 -435
rect 11388 -862 11393 -440
rect 11815 -862 11971 -440
rect 12393 -862 12399 -440
rect 11388 -867 11820 -862
rect -1320 -6240 -360 -6060
rect -1320 -6900 -1140 -6240
rect -480 -6900 -360 -6240
rect -1320 -9120 -360 -6900
rect -1320 -9900 -1140 -9120
rect -480 -9900 -360 -9120
rect -1320 -10140 -360 -9900
rect 2400 -6240 3360 -6060
rect 2400 -6900 2580 -6240
rect 3240 -6900 3360 -6240
rect 2400 -9120 3360 -6900
rect 2400 -9900 2580 -9120
rect 3240 -9900 3360 -9120
rect 2400 -10140 3360 -9900
rect -6054 -14352 -4864 -14150
rect -6054 -15078 -5790 -14352
rect -5098 -15078 -4864 -14352
rect -6054 -17042 -4864 -15078
rect -6054 -17966 -5794 -17042
rect -5118 -17966 -4864 -17042
rect -6054 -18246 -4864 -17966
<< via3 >>
rect 6352 16360 7028 17284
rect -1080 8460 -420 9240
rect 2640 8460 3300 9240
rect -8123 -112 -7797 214
rect 11971 -862 12393 -440
rect -1140 -9900 -480 -9120
rect 2580 -9900 3240 -9120
rect -5794 -17966 -5118 -17042
<< metal4 >>
rect 5418 24654 7998 25298
rect 5418 22976 5934 24654
rect 7354 22976 7998 24654
rect 5418 17284 7998 22976
rect 5418 16360 6352 17284
rect 7028 16360 7998 17284
rect 5418 15752 7998 16360
rect -1260 12660 -300 12900
rect -1260 12180 -1140 12660
rect -420 12180 -300 12660
rect -1260 9240 -300 12180
rect -1260 8460 -1080 9240
rect -420 8460 -300 9240
rect -1260 8100 -300 8460
rect 2460 12660 3420 12900
rect 2460 12180 2580 12660
rect 3300 12180 3420 12660
rect 2460 9240 3420 12180
rect 2460 8460 2640 9240
rect 3300 8460 3420 9240
rect 2460 8100 3420 8460
rect -8124 214 -7796 215
rect -8771 -112 -8123 214
rect -7797 -112 -7796 214
rect -8771 -391 -8445 -112
rect -8124 -113 -7796 -112
rect 11970 -440 12394 -439
rect 11970 -862 11971 -440
rect 12393 -862 13007 -440
rect 11970 -863 12394 -862
rect -1320 -9120 -360 -8760
rect -1320 -9900 -1140 -9120
rect -480 -9900 -360 -9120
rect -1320 -12840 -360 -9900
rect -1320 -13320 -1200 -12840
rect -480 -13320 -360 -12840
rect -1320 -13560 -360 -13320
rect 2400 -9120 3360 -8760
rect 2400 -9900 2580 -9120
rect 3240 -9900 3360 -9120
rect 2400 -12840 3360 -9900
rect 2400 -13320 2520 -12840
rect 3240 -13320 3360 -12840
rect 2400 -13560 3360 -13320
rect -6644 -17042 -4064 -16694
rect -6644 -17966 -5794 -17042
rect -5118 -17966 -4064 -17042
rect -6644 -23918 -4064 -17966
rect -6644 -25596 -6064 -23918
rect -4644 -25596 -4064 -23918
rect -6644 -26240 -4064 -25596
<< via4 >>
rect 5934 22976 7354 24654
rect -1140 12180 -420 12660
rect 2580 12180 3300 12660
rect -8771 -717 -8445 -391
rect 13007 -862 13429 -440
rect -1200 -13320 -480 -12840
rect 2520 -13320 3240 -12840
rect -6064 -25596 -4644 -23918
<< metal5 >>
rect -7104 25824 8896 42024
rect -28066 20160 -12066 25780
rect 5418 24654 7978 25824
rect 5418 22976 5934 24654
rect 7354 22976 7978 24654
rect 5418 22068 7978 22976
rect -28066 18900 -300 20160
rect 15120 20100 31120 25800
rect 14160 20084 31120 20100
rect 2392 18968 31120 20084
rect 2392 18952 5438 18968
rect 14160 18960 31120 18968
rect -28066 17000 -12066 18900
rect -28200 16000 -12060 17000
rect -28066 9580 -12066 16000
rect -1274 13080 -306 18900
rect -1294 12660 -284 13080
rect -1294 12180 -1140 12660
rect -420 12180 -284 12660
rect -1294 11980 -284 12180
rect 2426 12660 3436 18952
rect 2426 12180 2580 12660
rect 3300 12180 3436 12660
rect 2426 11980 3436 12180
rect 15120 9600 31120 18960
rect -28000 -86 -12000 7100
rect 15030 54 31030 7066
rect -28000 -391 -9774 -86
rect -8795 -391 -8421 -367
rect -28000 -717 -8771 -391
rect -8445 -717 -8421 -391
rect -28000 -1376 -9774 -717
rect -8795 -741 -8421 -717
rect 12734 -440 31030 54
rect 12734 -862 13007 -440
rect 13429 -862 31030 -440
rect -28000 -9100 -12000 -1376
rect 12734 -1486 31030 -862
rect 15030 -9134 31030 -1486
rect -28080 -19776 -12080 -11622
rect -1354 -12840 -344 -12640
rect -1354 -13320 -1200 -12840
rect -480 -13320 -344 -12840
rect -1354 -13740 -344 -13320
rect 2366 -12840 3376 -12640
rect 2366 -13320 2520 -12840
rect 3240 -13320 3376 -12840
rect -1334 -19776 -366 -13740
rect 2366 -19612 3376 -13320
rect 2332 -19628 5378 -19612
rect 15030 -19628 31030 -11764
rect -28080 -20702 -326 -19776
rect -28080 -27822 -12080 -20702
rect 2332 -20744 31030 -19628
rect 15002 -20852 31030 -20744
rect -6592 -23918 -4032 -23134
rect -6592 -25596 -6064 -23918
rect -4644 -25596 -4032 -23918
rect -6592 -27864 -4032 -25596
rect -7616 -44064 8384 -27864
rect 15030 -27964 31030 -20852
<< glass >>
rect -6800 26200 8600 41600
rect -27600 9800 -12466 25380
rect 15520 10000 30600 25400
rect -27600 -8700 -12400 6700
rect 15430 -8734 30630 6666
rect -27680 -27400 -12480 -12020
rect 15430 -27564 30630 -12164
rect -7200 -43800 8000 -28200
use GSense_nFET_6Contacts_V2  GSense_nFET_3VD_3Vg_5nf_V2_0
timestamp 1717352107
transform 1 0 315 0 1 -138
box 0 0 1 1
use GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH  GSense_nFET_3VD_3Vg_51nf_V2AllGates_VH_0
timestamp 1717386517
transform 1 0 -4684 0 1 542
box -1366 -1790 15678 80
<< end >>
