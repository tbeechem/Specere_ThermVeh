magic
tech sky130A
magscale 1 2
timestamp 1717301296
<< checkpaint >>
rect -1260 -1260 1267 1261
use not  x1
timestamp 0
transform 1 0 1 0 1 0
box 0 0 1 1
use not  x2
timestamp 0
transform 1 0 2 0 1 0
box 0 0 1 1
use not  x3
timestamp 0
transform 1 0 3 0 1 0
box 0 0 1 1
use not  x4
timestamp 0
transform 1 0 0 0 1 0
box 0 0 1 1
use not  x5
timestamp 0
transform 1 0 4 0 1 0
box 0 0 1 1
use not  x6
timestamp 0
transform 1 0 5 0 1 0
box 0 0 1 1
use not  x7
timestamp 0
transform 1 0 6 0 1 0
box 0 0 1 1
<< end >>
