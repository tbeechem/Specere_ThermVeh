magic
tech sky130A
magscale 1 2
timestamp 1717383051
<< pwell >>
rect 3214 -396 3295 -394
rect 3337 -396 3436 -382
rect 3214 -435 3436 -396
rect 3214 -485 3295 -435
rect 3337 -489 3436 -435
rect 13418 -484 13516 -202
rect 13688 -486 13786 -204
rect 3077 -696 3158 -665
rect 3077 -743 3251 -696
rect 3077 -744 3158 -743
<< locali >>
rect 162 -225 14659 -167
rect 161 -265 14659 -225
rect 161 -475 248 -265
rect 446 -476 544 -265
rect 722 -474 820 -265
rect 996 -478 1094 -265
rect 1274 -478 1372 -265
rect 1546 -476 1644 -265
rect 1824 -478 1922 -265
rect 2102 -478 2200 -265
rect 2380 -474 2478 -265
rect 2654 -478 2752 -265
rect 2930 -474 3028 -265
rect 3206 -474 3299 -455
rect 3484 -472 3582 -265
rect 3760 -482 3858 -265
rect 4032 -478 4130 -265
rect 4310 -478 4408 -265
rect 4582 -486 4680 -265
rect 4860 -478 4958 -265
rect 5136 -478 5234 -265
rect 5406 -480 5504 -265
rect 5692 -482 5790 -265
rect 5964 -482 6062 -265
rect 6244 -482 6342 -265
rect 6518 -482 6616 -265
rect 6794 -480 6892 -265
rect 7070 -482 7168 -265
rect 7346 -480 7444 -265
rect 7622 -480 7720 -265
rect 7898 -478 7996 -265
rect 8174 -480 8272 -265
rect 8450 -480 8548 -265
rect 8728 -480 8826 -265
rect 9004 -480 9102 -265
rect 9276 -482 9374 -265
rect 9554 -482 9652 -265
rect 9830 -478 9928 -265
rect 10108 -476 10206 -265
rect 10382 -480 10480 -265
rect 10658 -476 10756 -265
rect 10936 -476 11034 -265
rect 11212 -474 11310 -265
rect 11488 -478 11586 -265
rect 11764 -476 11862 -265
rect 12040 -476 12138 -265
rect 12314 -474 12412 -265
rect 12594 -474 12692 -265
rect 12870 -474 12968 -265
rect 13142 -474 13240 -265
rect 13418 -484 13516 -265
rect 13688 -486 13786 -265
rect 13980 -484 14078 -265
rect 169 -889 271 -649
rect 440 -889 538 -646
rect 712 -889 810 -650
rect 988 -889 1086 -654
rect 1266 -889 1364 -660
rect 1542 -889 1640 -664
rect 1816 -889 1914 -662
rect 2094 -889 2192 -664
rect 2372 -889 2470 -664
rect 2646 -889 2744 -664
rect 2924 -889 3022 -662
rect 3196 -692 3294 -654
rect 3472 -889 3570 -654
rect 3752 -889 3850 -660
rect 4020 -889 4118 -660
rect 4304 -889 4402 -664
rect 4578 -889 4676 -660
rect 4854 -889 4952 -664
rect 5128 -889 5226 -656
rect 5406 -889 5504 -664
rect 5676 -889 5774 -662
rect 5952 -889 6050 -656
rect 6234 -889 6332 -650
rect 6510 -889 6608 -654
rect 6784 -889 6882 -654
rect 7056 -889 7154 -654
rect 7338 -889 7436 -654
rect 7616 -889 7714 -660
rect 7890 -889 7988 -660
rect 8168 -889 8266 -664
rect 8444 -889 8542 -668
rect 8712 -889 8810 -668
rect 8994 -889 9092 -672
rect 9272 -889 9370 -670
rect 9546 -889 9644 -672
rect 9822 -889 9920 -672
rect 10092 -889 10190 -656
rect 10370 -889 10468 -664
rect 10652 -889 10750 -668
rect 10934 -889 11032 -664
rect 11202 -889 11300 -660
rect 11478 -889 11576 -660
rect 11748 -889 11846 -660
rect 12026 -889 12124 -654
rect 12308 -889 12406 -654
rect 12588 -889 12686 -654
rect 12854 -889 12952 -656
rect 13130 -889 13228 -662
rect 13410 -889 13508 -656
rect 13694 -889 13792 -656
rect 13972 -889 14070 -652
rect 14561 -889 14659 -265
rect 166 -920 14659 -889
rect 166 -976 4172 -920
rect 4250 -976 14659 -920
rect 166 -987 14659 -976
<< viali >>
rect 4172 -976 4250 -920
<< metal1 >>
rect 287 -348 15619 -282
rect -1366 -536 -1166 -400
rect -1366 -594 152 -536
rect -1366 -600 -1166 -594
rect -47 -772 -5 -594
rect 292 -614 332 -348
rect 374 -612 414 -348
rect 568 -772 598 -516
rect 654 -772 684 -516
rect 850 -612 890 -348
rect 918 -612 958 -348
rect 1122 -772 1152 -516
rect 1208 -772 1238 -516
rect 1398 -616 1438 -348
rect 1470 -612 1510 -348
rect 1670 -772 1700 -516
rect 1762 -772 1792 -518
rect 1950 -608 1990 -348
rect 2030 -608 2070 -348
rect 2220 -772 2250 -518
rect 2312 -772 2342 -520
rect 2504 -612 2544 -348
rect 2578 -610 2618 -348
rect 2776 -772 2806 -520
rect 2864 -772 2894 -522
rect 3056 -614 3096 -348
rect 3126 -610 3166 -348
rect 3337 -392 3436 -382
rect 3214 -396 3295 -394
rect 3337 -396 3352 -392
rect 3214 -435 3352 -396
rect 3214 -485 3295 -435
rect 3337 -472 3352 -435
rect 3426 -472 3436 -392
rect 3337 -489 3436 -472
rect 3211 -642 3285 -641
rect 3077 -677 3158 -665
rect 3077 -732 3088 -677
rect 3148 -696 3158 -677
rect 3200 -696 3291 -642
rect 3148 -732 3291 -696
rect 3077 -742 3291 -732
rect 3077 -743 3251 -742
rect 3077 -744 3158 -743
rect 3326 -772 3356 -522
rect 3414 -772 3444 -522
rect 3604 -614 3644 -348
rect 3682 -610 3722 -348
rect 3878 -772 3908 -520
rect 3966 -772 3996 -520
rect 4158 -622 4198 -348
rect 4236 -614 4276 -348
rect 4430 -772 4460 -520
rect 4522 -772 4552 -520
rect 4714 -612 4754 -348
rect 4788 -608 4828 -348
rect 4984 -772 5014 -510
rect 5070 -772 5100 -512
rect 5258 -612 5292 -348
rect 5348 -612 5382 -348
rect 5538 -772 5568 -514
rect 5624 -772 5654 -514
rect 5814 -612 5848 -348
rect 5898 -608 5932 -348
rect 6090 -772 6124 -510
rect 6172 -610 6206 -348
rect 6364 -772 6394 -512
rect 6452 -772 6482 -510
rect 6642 -608 6676 -348
rect 6728 -614 6762 -348
rect 6912 -772 6942 -510
rect 7004 -772 7034 -510
rect 7194 -606 7228 -348
rect 7280 -610 7314 -348
rect 7466 -772 7496 -510
rect 7558 -772 7588 -510
rect 7744 -610 7778 -348
rect 7832 -612 7866 -348
rect 8018 -772 8048 -510
rect 8104 -772 8134 -510
rect 8300 -616 8334 -348
rect 8382 -610 8416 -348
rect 8572 -772 8602 -510
rect 8660 -772 8690 -512
rect 8854 -612 8888 -348
rect 8932 -610 8966 -348
rect 9124 -772 9154 -508
rect 9212 -772 9242 -508
rect 9410 -620 9444 -348
rect 9484 -616 9518 -348
rect 9674 -772 9704 -506
rect 9762 -772 9792 -508
rect 9954 -620 9988 -348
rect 10034 -622 10068 -348
rect 10226 -772 10256 -508
rect 10314 -772 10344 -506
rect 10510 -620 10544 -348
rect 10584 -622 10618 -348
rect 10778 -772 10808 -508
rect 10868 -772 10898 -506
rect 11060 -618 11094 -348
rect 11136 -618 11170 -348
rect 11330 -772 11360 -508
rect 11420 -772 11450 -506
rect 11610 -614 11644 -348
rect 11692 -616 11726 -348
rect 11884 -772 11914 -502
rect 11974 -772 12004 -500
rect 12162 -610 12196 -348
rect 12240 -608 12274 -348
rect 12438 -772 12468 -500
rect 12524 -772 12554 -496
rect 12712 -612 12746 -348
rect 12796 -614 12830 -348
rect 12984 -772 13014 -510
rect 13076 -772 13106 -512
rect 13264 -612 13298 -348
rect 13348 -610 13382 -348
rect 13540 -772 13570 -510
rect 13624 -772 13654 -510
rect 13818 -606 13852 -348
rect 13896 -608 13930 -348
rect 14090 -772 14120 -510
rect 14210 -600 14244 -348
rect 15553 -474 15619 -348
rect 15478 -674 15678 -474
rect -47 -814 174 -772
rect 254 -814 14122 -772
rect 14080 -816 14122 -814
rect 4132 -920 4272 -908
rect 4132 -976 4172 -920
rect 4250 -976 4272 -920
rect 4132 -1590 4272 -976
rect 4118 -1790 4318 -1590
<< via1 >>
rect 3352 -472 3426 -392
rect 3088 -732 3148 -677
<< metal2 >>
rect 3264 404 3515 650
rect 3339 -392 3436 404
rect 3339 -472 3352 -392
rect 3426 -472 3436 -392
rect 3339 -491 3436 -472
rect 3077 -677 3159 -663
rect 3077 -732 3088 -677
rect 3148 -732 3159 -677
rect 3077 -1578 3159 -732
rect 2970 -1793 3189 -1578
rect 3077 -1797 3159 -1793
use sky130_fd_pr__nfet_03v3_nvt_XW2EXC  XM1 ~/Specere_ThermVeh/mag
timestamp 1717383051
transform 1 0 7113 0 1 -566
box -7178 -300 7178 300
<< labels >>
flabel metal1 4118 -1790 4318 -1590 0 FreeSans 256 0 0 0 VG_H
port 0 nsew
flabel metal1 -1366 -600 -1166 -400 0 FreeSans 256 0 0 0 VD_H
port 1 nsew
flabel metal1 15478 -674 15678 -474 0 FreeSans 256 0 0 0 VLow_Src
port 2 nsew
<< end >>
